
`ifndef IDI_NUM
    `define IDI_NUM 4
`endif

`ifndef AGG_NUM
    `define AGG_NUM 4
`endif

`define AGG_PATH as6d_app_tb.u_as6d_app
