
`include "as6d_app_all_includes.vh"
//`include "as6d_mep_all_includes.vh"
module   as6d_app_video_pipe #(
	parameter	VIDEO_DATA_SIZE		= 140,
	parameter	DATA_PARITY_WIDTH	= 21
)(/*AUTOARG*/
   // Outputs
   video_pipe_date_type_for_concat_align_vld7,
   video_pipe_date_type_for_concat_align_vld6,
   video_pipe_date_type_for_concat_align_vld5,
   video_pipe_date_type_for_concat_align_vld4,
   video_pipe_date_type_for_concat_align_vld3,
   video_pipe_date_type_for_concat_align_vld2,
   video_pipe_date_type_for_concat_align_vld1,
   video_pipe_date_type_for_concat_align_vld0,
   video_pipe_date_type_for_concat_align7,
   video_pipe_date_type_for_concat_align6,
   video_pipe_date_type_for_concat_align5,
   video_pipe_date_type_for_concat_align4,
   video_pipe_date_type_for_concat_align3,
   video_pipe_date_type_for_concat_align2,
   video_pipe_date_type_for_concat_align1,
   video_pipe_date_type_for_concat_align0,
   video_pipe7_vld_aggre_bypass, video_pipe7_data_aggre_bypass,
   video_pipe6_vld_aggre_bypass, video_pipe6_data_aggre_bypass,
   video_pipe5_vld_aggre_bypass, video_pipe5_data_aggre_bypass,
   video_pipe4_vld_aggre_bypass, video_pipe4_data_aggre_bypass,
   video_pipe3_vld_aggre_bypass, video_pipe3_data_aggre_bypass,
   video_pipe2_vld_aggre_bypass, video_pipe2_data_aggre_bypass,
   video_pipe1_vld_aggre_bypass, video_pipe1_data_aggre_bypass,
   video_pipe0_vld_aggre_bypass, video_pipe0_data_aggre_bypass,
   video_loss7, video_loss6, video_loss5, video_loss4, video_loss3,
   video_loss2, video_loss1, video_loss0, video_lock7, video_lock6,
   video_lock5, video_lock4, video_lock3, video_lock2, video_lock1,
   video_lock0, video_data_vld7, video_data_vld6, video_data_vld5,
   video_data_vld4, video_data_vld3, video_data_vld2, video_data_vld1,
   video_data_vld0, video_data_fwft_fifo_udf_int7,
   video_data_fwft_fifo_udf_int6, video_data_fwft_fifo_udf_int5,
   video_data_fwft_fifo_udf_int4, video_data_fwft_fifo_udf_int3,
   video_data_fwft_fifo_udf_int2, video_data_fwft_fifo_udf_int1,
   video_data_fwft_fifo_udf_int0, video_data_fwft_fifo_single_err7,
   video_data_fwft_fifo_single_err6, video_data_fwft_fifo_single_err5,
   video_data_fwft_fifo_single_err4, video_data_fwft_fifo_single_err3,
   video_data_fwft_fifo_single_err2, video_data_fwft_fifo_single_err1,
   video_data_fwft_fifo_single_err0, video_data_fwft_fifo_prog_full7,
   video_data_fwft_fifo_prog_full6, video_data_fwft_fifo_prog_full5,
   video_data_fwft_fifo_prog_full4, video_data_fwft_fifo_prog_full3,
   video_data_fwft_fifo_prog_full2, video_data_fwft_fifo_prog_full1,
   video_data_fwft_fifo_prog_full0, video_data_fwft_fifo_ovf_int7,
   video_data_fwft_fifo_ovf_int6, video_data_fwft_fifo_ovf_int5,
   video_data_fwft_fifo_ovf_int4, video_data_fwft_fifo_ovf_int3,
   video_data_fwft_fifo_ovf_int2, video_data_fwft_fifo_ovf_int1,
   video_data_fwft_fifo_ovf_int0, video_data_fwft_fifo_full7,
   video_data_fwft_fifo_full6, video_data_fwft_fifo_full5,
   video_data_fwft_fifo_full4, video_data_fwft_fifo_full3,
   video_data_fwft_fifo_full2, video_data_fwft_fifo_full1,
   video_data_fwft_fifo_full0, video_data_fwft_fifo_empty7,
   video_data_fwft_fifo_empty6, video_data_fwft_fifo_empty5,
   video_data_fwft_fifo_empty4, video_data_fwft_fifo_empty3,
   video_data_fwft_fifo_empty2, video_data_fwft_fifo_empty1,
   video_data_fwft_fifo_empty0, video_data_fwft_fifo_ecc_fault7,
   video_data_fwft_fifo_ecc_fault6, video_data_fwft_fifo_ecc_fault5,
   video_data_fwft_fifo_ecc_fault4, video_data_fwft_fifo_ecc_fault3,
   video_data_fwft_fifo_ecc_fault2, video_data_fwft_fifo_ecc_fault1,
   video_data_fwft_fifo_ecc_fault0, video_data_fwft_fifo_double_err7,
   video_data_fwft_fifo_double_err6, video_data_fwft_fifo_double_err5,
   video_data_fwft_fifo_double_err4, video_data_fwft_fifo_double_err3,
   video_data_fwft_fifo_double_err2, video_data_fwft_fifo_double_err1,
   video_data_fwft_fifo_double_err0, video_data_afifo_udf_int7,
   video_data_afifo_udf_int6, video_data_afifo_udf_int5,
   video_data_afifo_udf_int4, video_data_afifo_udf_int3,
   video_data_afifo_udf_int2, video_data_afifo_udf_int1,
   video_data_afifo_udf_int0, video_data_afifo_single_err7,
   video_data_afifo_single_err6, video_data_afifo_single_err5,
   video_data_afifo_single_err4, video_data_afifo_single_err3,
   video_data_afifo_single_err2, video_data_afifo_single_err1,
   video_data_afifo_single_err0, video_data_afifo_prog_full7,
   video_data_afifo_prog_full6, video_data_afifo_prog_full5,
   video_data_afifo_prog_full4, video_data_afifo_prog_full3,
   video_data_afifo_prog_full2, video_data_afifo_prog_full1,
   video_data_afifo_prog_full0, video_data_afifo_prog_empty7,
   video_data_afifo_prog_empty6, video_data_afifo_prog_empty5,
   video_data_afifo_prog_empty4, video_data_afifo_prog_empty3,
   video_data_afifo_prog_empty2, video_data_afifo_prog_empty1,
   video_data_afifo_prog_empty0, video_data_afifo_ovf_int7,
   video_data_afifo_ovf_int6, video_data_afifo_ovf_int5,
   video_data_afifo_ovf_int4, video_data_afifo_ovf_int3,
   video_data_afifo_ovf_int2, video_data_afifo_ovf_int1,
   video_data_afifo_ovf_int0, video_data_afifo_full7,
   video_data_afifo_full6, video_data_afifo_full5,
   video_data_afifo_full4, video_data_afifo_full3,
   video_data_afifo_full2, video_data_afifo_full1,
   video_data_afifo_full0, video_data_afifo_empty7,
   video_data_afifo_empty6, video_data_afifo_empty5,
   video_data_afifo_empty4, video_data_afifo_empty3,
   video_data_afifo_empty2, video_data_afifo_empty1,
   video_data_afifo_empty0, video_data_afifo_ecc_fault7,
   video_data_afifo_ecc_fault6, video_data_afifo_ecc_fault5,
   video_data_afifo_ecc_fault4, video_data_afifo_ecc_fault3,
   video_data_afifo_ecc_fault2, video_data_afifo_ecc_fault1,
   video_data_afifo_ecc_fault0, video_data_afifo_double_err7,
   video_data_afifo_double_err6, video_data_afifo_double_err5,
   video_data_afifo_double_err4, video_data_afifo_double_err3,
   video_data_afifo_double_err2, video_data_afifo_double_err1,
   video_data_afifo_double_err0, video_data7, video_data6,
   video_data5, video_data4, video_data3, video_data2, video_data1,
   video_data0, reg_rd_resv_pkt_cnt_sp_ls_pipe7,
   reg_rd_resv_pkt_cnt_sp_ls_pipe6, reg_rd_resv_pkt_cnt_sp_ls_pipe5,
   reg_rd_resv_pkt_cnt_sp_ls_pipe4, reg_rd_resv_pkt_cnt_sp_ls_pipe3,
   reg_rd_resv_pkt_cnt_sp_ls_pipe2, reg_rd_resv_pkt_cnt_sp_ls_pipe1,
   reg_rd_resv_pkt_cnt_sp_ls_pipe0, reg_rd_resv_pkt_cnt_sp_le_pipe7,
   reg_rd_resv_pkt_cnt_sp_le_pipe6, reg_rd_resv_pkt_cnt_sp_le_pipe5,
   reg_rd_resv_pkt_cnt_sp_le_pipe4, reg_rd_resv_pkt_cnt_sp_le_pipe3,
   reg_rd_resv_pkt_cnt_sp_le_pipe2, reg_rd_resv_pkt_cnt_sp_le_pipe1,
   reg_rd_resv_pkt_cnt_sp_le_pipe0, reg_rd_resv_pkt_cnt_sp_fs_pipe7,
   reg_rd_resv_pkt_cnt_sp_fs_pipe6, reg_rd_resv_pkt_cnt_sp_fs_pipe5,
   reg_rd_resv_pkt_cnt_sp_fs_pipe4, reg_rd_resv_pkt_cnt_sp_fs_pipe3,
   reg_rd_resv_pkt_cnt_sp_fs_pipe2, reg_rd_resv_pkt_cnt_sp_fs_pipe1,
   reg_rd_resv_pkt_cnt_sp_fs_pipe0, reg_rd_resv_pkt_cnt_sp_fe_pipe7,
   reg_rd_resv_pkt_cnt_sp_fe_pipe6, reg_rd_resv_pkt_cnt_sp_fe_pipe5,
   reg_rd_resv_pkt_cnt_sp_fe_pipe4, reg_rd_resv_pkt_cnt_sp_fe_pipe3,
   reg_rd_resv_pkt_cnt_sp_fe_pipe2, reg_rd_resv_pkt_cnt_sp_fe_pipe1,
   reg_rd_resv_pkt_cnt_sp_fe_pipe0, reg_rd_resv_pkt_cnt_lp_ph_pipe7,
   reg_rd_resv_pkt_cnt_lp_ph_pipe6, reg_rd_resv_pkt_cnt_lp_ph_pipe5,
   reg_rd_resv_pkt_cnt_lp_ph_pipe4, reg_rd_resv_pkt_cnt_lp_ph_pipe3,
   reg_rd_resv_pkt_cnt_lp_ph_pipe2, reg_rd_resv_pkt_cnt_lp_ph_pipe1,
   reg_rd_resv_pkt_cnt_lp_ph_pipe0, reg_rd_resv_pkt_cnt_lp_pf_pipe7,
   reg_rd_resv_pkt_cnt_lp_pf_pipe6, reg_rd_resv_pkt_cnt_lp_pf_pipe5,
   reg_rd_resv_pkt_cnt_lp_pf_pipe4, reg_rd_resv_pkt_cnt_lp_pf_pipe3,
   reg_rd_resv_pkt_cnt_lp_pf_pipe2, reg_rd_resv_pkt_cnt_lp_pf_pipe1,
   reg_rd_resv_pkt_cnt_lp_pf_pipe0,
   reg_rd_pipe7_dispatched_cnt_ready_for_sch,
   reg_rd_pipe6_dispatched_cnt_ready_for_sch,
   reg_rd_pipe5_dispatched_cnt_ready_for_sch,
   reg_rd_pipe4_dispatched_cnt_ready_for_sch,
   reg_rd_pipe3_dispatched_cnt_ready_for_sch,
   reg_rd_pipe2_dispatched_cnt_ready_for_sch,
   reg_rd_pipe1_dispatched_cnt_ready_for_sch,
   reg_rd_pipe0_dispatched_cnt_ready_for_sch,
   reg_rd_dbg_pkt_num_nonzero_threshold_err,
   reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err,
   reg_rd_app_full_cnt_sync_fifo_pipe7,
   reg_rd_app_full_cnt_sync_fifo_pipe6,
   reg_rd_app_full_cnt_sync_fifo_pipe5,
   reg_rd_app_full_cnt_sync_fifo_pipe4,
   reg_rd_app_full_cnt_sync_fifo_pipe3,
   reg_rd_app_full_cnt_sync_fifo_pipe2,
   reg_rd_app_full_cnt_sync_fifo_pipe1,
   reg_rd_app_full_cnt_sync_fifo_pipe0,
   reg_rd_app_full_cnt_async_fifo_pipe7,
   reg_rd_app_full_cnt_async_fifo_pipe6,
   reg_rd_app_full_cnt_async_fifo_pipe5,
   reg_rd_app_full_cnt_async_fifo_pipe4,
   reg_rd_app_full_cnt_async_fifo_pipe3,
   reg_rd_app_full_cnt_async_fifo_pipe2,
   reg_rd_app_full_cnt_async_fifo_pipe1,
   reg_rd_app_full_cnt_async_fifo_pipe0,
   line_end_vld_pipe7_aggregator3, line_end_vld_pipe7_aggregator2,
   line_end_vld_pipe7_aggregator1, line_end_vld_pipe7_aggregator0,
   line_end_vld_pipe6_aggregator3, line_end_vld_pipe6_aggregator2,
   line_end_vld_pipe6_aggregator1, line_end_vld_pipe6_aggregator0,
   line_end_vld_pipe5_aggregator3, line_end_vld_pipe5_aggregator2,
   line_end_vld_pipe5_aggregator1, line_end_vld_pipe5_aggregator0,
   line_end_vld_pipe4_aggregator3, line_end_vld_pipe4_aggregator2,
   line_end_vld_pipe4_aggregator1, line_end_vld_pipe4_aggregator0,
   line_end_vld_pipe3_aggregator3, line_end_vld_pipe3_aggregator2,
   line_end_vld_pipe3_aggregator1, line_end_vld_pipe3_aggregator0,
   line_end_vld_pipe2_aggregator3, line_end_vld_pipe2_aggregator2,
   line_end_vld_pipe2_aggregator1, line_end_vld_pipe2_aggregator0,
   line_end_vld_pipe1_aggregator3, line_end_vld_pipe1_aggregator2,
   line_end_vld_pipe1_aggregator1, line_end_vld_pipe1_aggregator0,
   line_end_vld_pipe0_aggregator3, line_end_vld_pipe0_aggregator2,
   line_end_vld_pipe0_aggregator1, line_end_vld_pipe0_aggregator0,
   line_end7, line_end6, line_end5, line_end4, line_end3, line_end2,
   line_end1, line_end0, lcrc_err7, lcrc_err6, lcrc_err5, lcrc_err4,
   lcrc_err3, lcrc_err2, lcrc_err1, lcrc_err0, fs_detect_pipe7,
   fs_detect_pipe6, fs_detect_pipe5, fs_detect_pipe4, fs_detect_pipe3,
   fs_detect_pipe2, fs_detect_pipe1, fs_detect_pipe0, fs_cnt_pipe7,
   fs_cnt_pipe6, fs_cnt_pipe5, fs_cnt_pipe4, fs_cnt_pipe3,
   fs_cnt_pipe2, fs_cnt_pipe1, fs_cnt_pipe0, fifo_rd_ctrl_cs7,
   fifo_rd_ctrl_cs6, fifo_rd_ctrl_cs5, fifo_rd_ctrl_cs4,
   fifo_rd_ctrl_cs3, fifo_rd_ctrl_cs2, fifo_rd_ctrl_cs1,
   fifo_rd_ctrl_cs0, empty_vld_pipe7_aggregator3,
   empty_vld_pipe7_aggregator2, empty_vld_pipe7_aggregator1,
   empty_vld_pipe7_aggregator0, empty_vld_pipe6_aggregator3,
   empty_vld_pipe6_aggregator2, empty_vld_pipe6_aggregator1,
   empty_vld_pipe6_aggregator0, empty_vld_pipe5_aggregator3,
   empty_vld_pipe5_aggregator2, empty_vld_pipe5_aggregator1,
   empty_vld_pipe5_aggregator0, empty_vld_pipe4_aggregator3,
   empty_vld_pipe4_aggregator2, empty_vld_pipe4_aggregator1,
   empty_vld_pipe4_aggregator0, empty_vld_pipe3_aggregator3,
   empty_vld_pipe3_aggregator2, empty_vld_pipe3_aggregator1,
   empty_vld_pipe3_aggregator0, empty_vld_pipe2_aggregator3,
   empty_vld_pipe2_aggregator2, empty_vld_pipe2_aggregator1,
   empty_vld_pipe2_aggregator0, empty_vld_pipe1_aggregator3,
   empty_vld_pipe1_aggregator2, empty_vld_pipe1_aggregator1,
   empty_vld_pipe1_aggregator0, empty_vld_pipe0_aggregator3,
   empty_vld_pipe0_aggregator2, empty_vld_pipe0_aggregator1,
   empty_vld_pipe0_aggregator0, ack_vld_pipe7_aggregator3,
   ack_vld_pipe7_aggregator2, ack_vld_pipe7_aggregator1,
   ack_vld_pipe7_aggregator0, ack_vld_pipe6_aggregator3,
   ack_vld_pipe6_aggregator2, ack_vld_pipe6_aggregator1,
   ack_vld_pipe6_aggregator0, ack_vld_pipe5_aggregator3,
   ack_vld_pipe5_aggregator2, ack_vld_pipe5_aggregator1,
   ack_vld_pipe5_aggregator0, ack_vld_pipe4_aggregator3,
   ack_vld_pipe4_aggregator2, ack_vld_pipe4_aggregator1,
   ack_vld_pipe4_aggregator0, ack_vld_pipe3_aggregator3,
   ack_vld_pipe3_aggregator2, ack_vld_pipe3_aggregator1,
   ack_vld_pipe3_aggregator0, ack_vld_pipe2_aggregator3,
   ack_vld_pipe2_aggregator2, ack_vld_pipe2_aggregator1,
   ack_vld_pipe2_aggregator0, ack_vld_pipe1_aggregator3,
   ack_vld_pipe1_aggregator2, ack_vld_pipe1_aggregator1,
   ack_vld_pipe1_aggregator0, ack_vld_pipe0_aggregator3,
   ack_vld_pipe0_aggregator2, ack_vld_pipe0_aggregator1,
   ack_vld_pipe0_aggregator0, ack_pre7, ack_pre6, ack_pre5, ack_pre4,
   ack_pre3, ack_pre2, ack_pre1, ack_pre0, ack7, ack6, ack5, ack4,
   ack3, ack2, ack1, ack0, reg_rd_pipe_fifo_full,
   // Inputs
   video_loss_en7, video_loss_en6, video_loss_en5, video_loss_en4,
   video_loss_en3, video_loss_en2, video_loss_en1, video_loss_en0,
   up_state_video_pipe7, up_state_video_pipe6, up_state_video_pipe5,
   up_state_video_pipe4, up_state_video_pipe3, up_state_video_pipe2,
   up_state_video_pipe1, up_state_video_pipe0, time_window7,
   time_window6, time_window5, time_window4, time_window3,
   time_window2, time_window1, time_window0, reg_video_pipe_en,
   reg_video_fifo_empty_depend_cnt_mux, reg_sram_lcrc_err_oen,
   reg_resv_pkt_match_lp_dt_pipe7, reg_resv_pkt_match_lp_dt_pipe6,
   reg_resv_pkt_match_lp_dt_pipe5, reg_resv_pkt_match_lp_dt_pipe4,
   reg_resv_pkt_match_lp_dt_pipe3, reg_resv_pkt_match_lp_dt_pipe2,
   reg_resv_pkt_match_lp_dt_pipe1, reg_resv_pkt_match_lp_dt_pipe0,
   reg_resv_pkt_match_lp_dt_en_pipe7,
   reg_resv_pkt_match_lp_dt_en_pipe6,
   reg_resv_pkt_match_lp_dt_en_pipe5,
   reg_resv_pkt_match_lp_dt_en_pipe4,
   reg_resv_pkt_match_lp_dt_en_pipe3,
   reg_resv_pkt_match_lp_dt_en_pipe2,
   reg_resv_pkt_match_lp_dt_en_pipe1,
   reg_resv_pkt_match_lp_dt_en_pipe0, reg_last_byte_header_down_mux,
   reg_dft_tpram_config, reg_dft_sync_tpram_config,
   reg_dbg_pkt_num_nonzero_threshold,
   reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold,
   reg_clear_resv_pkt_cnt_sp_ls_pipe7,
   reg_clear_resv_pkt_cnt_sp_ls_pipe6,
   reg_clear_resv_pkt_cnt_sp_ls_pipe5,
   reg_clear_resv_pkt_cnt_sp_ls_pipe4,
   reg_clear_resv_pkt_cnt_sp_ls_pipe3,
   reg_clear_resv_pkt_cnt_sp_ls_pipe2,
   reg_clear_resv_pkt_cnt_sp_ls_pipe1,
   reg_clear_resv_pkt_cnt_sp_ls_pipe0,
   reg_clear_resv_pkt_cnt_sp_le_pipe7,
   reg_clear_resv_pkt_cnt_sp_le_pipe6,
   reg_clear_resv_pkt_cnt_sp_le_pipe5,
   reg_clear_resv_pkt_cnt_sp_le_pipe4,
   reg_clear_resv_pkt_cnt_sp_le_pipe3,
   reg_clear_resv_pkt_cnt_sp_le_pipe2,
   reg_clear_resv_pkt_cnt_sp_le_pipe1,
   reg_clear_resv_pkt_cnt_sp_le_pipe0,
   reg_clear_resv_pkt_cnt_sp_fs_pipe7,
   reg_clear_resv_pkt_cnt_sp_fs_pipe6,
   reg_clear_resv_pkt_cnt_sp_fs_pipe5,
   reg_clear_resv_pkt_cnt_sp_fs_pipe4,
   reg_clear_resv_pkt_cnt_sp_fs_pipe3,
   reg_clear_resv_pkt_cnt_sp_fs_pipe2,
   reg_clear_resv_pkt_cnt_sp_fs_pipe1,
   reg_clear_resv_pkt_cnt_sp_fs_pipe0,
   reg_clear_resv_pkt_cnt_sp_fe_pipe7,
   reg_clear_resv_pkt_cnt_sp_fe_pipe6,
   reg_clear_resv_pkt_cnt_sp_fe_pipe5,
   reg_clear_resv_pkt_cnt_sp_fe_pipe4,
   reg_clear_resv_pkt_cnt_sp_fe_pipe3,
   reg_clear_resv_pkt_cnt_sp_fe_pipe2,
   reg_clear_resv_pkt_cnt_sp_fe_pipe1,
   reg_clear_resv_pkt_cnt_sp_fe_pipe0,
   reg_clear_resv_pkt_cnt_lp_ph_pipe7,
   reg_clear_resv_pkt_cnt_lp_ph_pipe6,
   reg_clear_resv_pkt_cnt_lp_ph_pipe5,
   reg_clear_resv_pkt_cnt_lp_ph_pipe4,
   reg_clear_resv_pkt_cnt_lp_ph_pipe3,
   reg_clear_resv_pkt_cnt_lp_ph_pipe2,
   reg_clear_resv_pkt_cnt_lp_ph_pipe1,
   reg_clear_resv_pkt_cnt_lp_ph_pipe0,
   reg_clear_resv_pkt_cnt_lp_pf_pipe7,
   reg_clear_resv_pkt_cnt_lp_pf_pipe6,
   reg_clear_resv_pkt_cnt_lp_pf_pipe5,
   reg_clear_resv_pkt_cnt_lp_pf_pipe4,
   reg_clear_resv_pkt_cnt_lp_pf_pipe3,
   reg_clear_resv_pkt_cnt_lp_pf_pipe2,
   reg_clear_resv_pkt_cnt_lp_pf_pipe1,
   reg_clear_resv_pkt_cnt_lp_pf_pipe0,
   reg_clear_app_full_cnt_sync_fifo_pipe7,
   reg_clear_app_full_cnt_sync_fifo_pipe6,
   reg_clear_app_full_cnt_sync_fifo_pipe5,
   reg_clear_app_full_cnt_sync_fifo_pipe4,
   reg_clear_app_full_cnt_sync_fifo_pipe3,
   reg_clear_app_full_cnt_sync_fifo_pipe2,
   reg_clear_app_full_cnt_sync_fifo_pipe1,
   reg_clear_app_full_cnt_sync_fifo_pipe0,
   reg_clear_app_full_cnt_async_fifo_pipe7,
   reg_clear_app_full_cnt_async_fifo_pipe6,
   reg_clear_app_full_cnt_async_fifo_pipe5,
   reg_clear_app_full_cnt_async_fifo_pipe4,
   reg_clear_app_full_cnt_async_fifo_pipe3,
   reg_clear_app_full_cnt_async_fifo_pipe2,
   reg_clear_app_full_cnt_async_fifo_pipe1,
   reg_clear_app_full_cnt_async_fifo_pipe0,
   reg_app_wr_idi_data_continue, reg_app_pkt_crc_gen_dis,
   reg_app_ecc_fault_detc_en, reg_app_ecc_bypass,
   reg_app_ecc_addr_protect_en, pipe7_word_count,
   pipe7_virtual_channel_x, pipe7_virtual_channel, pipe7_pkt_crc_en,
   pipe7_pkt_crc, pipe7_header_en, pipe7_data_type, pipe7_data_en,
   pipe7_csi_data, pipe7_bytes_en, pipe7_aggr_id, pipe6_word_count,
   pipe6_virtual_channel_x, pipe6_virtual_channel, pipe6_pkt_crc_en,
   pipe6_pkt_crc, pipe6_header_en, pipe6_data_type, pipe6_data_en,
   pipe6_csi_data, pipe6_bytes_en, pipe6_aggr_id, pipe5_word_count,
   pipe5_virtual_channel_x, pipe5_virtual_channel, pipe5_pkt_crc_en,
   pipe5_pkt_crc, pipe5_header_en, pipe5_data_type, pipe5_data_en,
   pipe5_csi_data, pipe5_bytes_en, pipe5_aggr_id, pipe4_word_count,
   pipe4_virtual_channel_x, pipe4_virtual_channel, pipe4_pkt_crc_en,
   pipe4_pkt_crc, pipe4_header_en, pipe4_data_type, pipe4_data_en,
   pipe4_csi_data, pipe4_bytes_en, pipe4_aggr_id, pipe3_word_count,
   pipe3_virtual_channel_x, pipe3_virtual_channel, pipe3_pkt_crc_en,
   pipe3_pkt_crc, pipe3_header_en, pipe3_data_type, pipe3_data_en,
   pipe3_csi_data, pipe3_bytes_en, pipe3_aggr_id, pipe2_word_count,
   pipe2_virtual_channel_x, pipe2_virtual_channel, pipe2_pkt_crc_en,
   pipe2_pkt_crc, pipe2_header_en, pipe2_data_type, pipe2_data_en,
   pipe2_csi_data, pipe2_bytes_en, pipe2_aggr_id, pipe1_word_count,
   pipe1_virtual_channel_x, pipe1_virtual_channel, pipe1_pkt_crc_en,
   pipe1_pkt_crc, pipe1_header_en, pipe1_data_type, pipe1_data_en,
   pipe1_csi_data, pipe1_bytes_en, pipe1_aggr_id, pipe0_word_count,
   pipe0_virtual_channel_x, pipe0_virtual_channel, pipe0_pkt_crc_en,
   pipe0_pkt_crc, pipe0_header_en, pipe0_data_type, pipe0_data_en,
   pipe0_csi_data, pipe0_bytes_en, pipe0_aggr_id, line_delay_en7,
   line_delay_en6, line_delay_en5, line_delay_en4, line_delay_en3,
   line_delay_en2, line_delay_en1, line_delay_en0, fifo_wrclk_rst_n7,
   fifo_wrclk_rst_n6, fifo_wrclk_rst_n5, fifo_wrclk_rst_n4,
   fifo_wrclk_rst_n3, fifo_wrclk_rst_n2, fifo_wrclk_rst_n1,
   fifo_wrclk_rst_n0, fifo_wrclk7, fifo_wrclk6, fifo_wrclk5,
   fifo_wrclk4, fifo_wrclk3, fifo_wrclk2, fifo_wrclk1, fifo_wrclk0,
   fifo_rdclk_rst_n7, fifo_rdclk_rst_n6, fifo_rdclk_rst_n5,
   fifo_rdclk_rst_n4, fifo_rdclk_rst_n3, fifo_rdclk_rst_n2,
   fifo_rdclk_rst_n1, fifo_rdclk_rst_n0, fifo_rdclk7, fifo_rdclk6,
   fifo_rdclk5, fifo_rdclk4, fifo_rdclk3, fifo_rdclk2, fifo_rdclk1,
   fifo_rdclk0, clk_1M, app_aggregation_bypass, pipe_fifo_full_clear
   );


/*AUTOINPUT*/
// Beginning of automatic inputs (from unused autoinst inputs)
input			app_aggregation_bypass;	// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input			clk_1M;			// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input			fifo_rdclk0;		// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk1;		// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk2;		// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk3;		// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk4;		// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk5;		// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk6;		// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk7;		// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk_rst_n0;	// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk_rst_n1;	// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk_rst_n2;	// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk_rst_n3;	// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk_rst_n4;	// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk_rst_n5;	// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk_rst_n6;	// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_rdclk_rst_n7;	// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk0;		// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk1;		// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk2;		// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk3;		// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk4;		// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk5;		// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk6;		// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk7;		// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk_rst_n0;	// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk_rst_n1;	// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk_rst_n2;	// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk_rst_n3;	// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk_rst_n4;	// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk_rst_n5;	// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk_rst_n6;	// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			fifo_wrclk_rst_n7;	// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			line_delay_en0;		// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			line_delay_en1;		// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			line_delay_en2;		// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			line_delay_en3;		// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			line_delay_en4;		// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			line_delay_en5;		// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			line_delay_en6;		// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			line_delay_en7;		// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [3:0]		pipe0_aggr_id;		// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0] pipe0_bytes_en;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0] pipe0_csi_data;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe0_data_en;		// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		pipe0_data_type;	// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe0_header_en;	// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [31:0]		pipe0_pkt_crc;		// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe0_pkt_crc_en;	// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [1:0]		pipe0_virtual_channel;	// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0] pipe0_virtual_channel_x;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [15:0]		pipe0_word_count;	// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [3:0]		pipe1_aggr_id;		// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0] pipe1_bytes_en;// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0] pipe1_csi_data;// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe1_data_en;		// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		pipe1_data_type;	// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe1_header_en;	// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [31:0]		pipe1_pkt_crc;		// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe1_pkt_crc_en;	// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [1:0]		pipe1_virtual_channel;	// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0] pipe1_virtual_channel_x;// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [15:0]		pipe1_word_count;	// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [3:0]		pipe2_aggr_id;		// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0] pipe2_bytes_en;// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0] pipe2_csi_data;// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe2_data_en;		// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		pipe2_data_type;	// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe2_header_en;	// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [31:0]		pipe2_pkt_crc;		// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe2_pkt_crc_en;	// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [1:0]		pipe2_virtual_channel;	// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0] pipe2_virtual_channel_x;// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [15:0]		pipe2_word_count;	// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [3:0]		pipe3_aggr_id;		// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0] pipe3_bytes_en;// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0] pipe3_csi_data;// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe3_data_en;		// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		pipe3_data_type;	// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe3_header_en;	// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [31:0]		pipe3_pkt_crc;		// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe3_pkt_crc_en;	// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [1:0]		pipe3_virtual_channel;	// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0] pipe3_virtual_channel_x;// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [15:0]		pipe3_word_count;	// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [3:0]		pipe4_aggr_id;		// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0] pipe4_bytes_en;// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0] pipe4_csi_data;// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe4_data_en;		// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		pipe4_data_type;	// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe4_header_en;	// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [31:0]		pipe4_pkt_crc;		// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe4_pkt_crc_en;	// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [1:0]		pipe4_virtual_channel;	// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0] pipe4_virtual_channel_x;// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [15:0]		pipe4_word_count;	// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [3:0]		pipe5_aggr_id;		// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0] pipe5_bytes_en;// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0] pipe5_csi_data;// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe5_data_en;		// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		pipe5_data_type;	// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe5_header_en;	// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [31:0]		pipe5_pkt_crc;		// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe5_pkt_crc_en;	// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [1:0]		pipe5_virtual_channel;	// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0] pipe5_virtual_channel_x;// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [15:0]		pipe5_word_count;	// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [3:0]		pipe6_aggr_id;		// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0] pipe6_bytes_en;// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0] pipe6_csi_data;// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe6_data_en;		// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		pipe6_data_type;	// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe6_header_en;	// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [31:0]		pipe6_pkt_crc;		// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe6_pkt_crc_en;	// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [1:0]		pipe6_virtual_channel;	// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0] pipe6_virtual_channel_x;// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [15:0]		pipe6_word_count;	// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [3:0]		pipe7_aggr_id;		// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0] pipe7_bytes_en;// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0] pipe7_csi_data;// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe7_data_en;		// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		pipe7_data_type;	// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe7_header_en;	// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [31:0]		pipe7_pkt_crc;		// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			pipe7_pkt_crc_en;	// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [1:0]		pipe7_virtual_channel;	// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0] pipe7_virtual_channel_x;// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [15:0]		pipe7_word_count;	// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_app_ecc_addr_protect_en;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input			reg_app_ecc_bypass;	// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input			reg_app_ecc_fault_detc_en;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input			reg_app_pkt_crc_gen_dis;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input			reg_app_wr_idi_data_continue;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input			reg_clear_app_full_cnt_async_fifo_pipe0;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_async_fifo_pipe1;// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_async_fifo_pipe2;// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_async_fifo_pipe3;// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_async_fifo_pipe4;// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_async_fifo_pipe5;// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_async_fifo_pipe6;// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_async_fifo_pipe7;// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_sync_fifo_pipe0;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_sync_fifo_pipe1;// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_sync_fifo_pipe2;// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_sync_fifo_pipe3;// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_sync_fifo_pipe4;// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_sync_fifo_pipe5;// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_sync_fifo_pipe6;// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_app_full_cnt_sync_fifo_pipe7;// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_pf_pipe0;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_pf_pipe1;// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_pf_pipe2;// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_pf_pipe3;// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_pf_pipe4;// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_pf_pipe5;// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_pf_pipe6;// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_pf_pipe7;// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_ph_pipe0;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_ph_pipe1;// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_ph_pipe2;// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_ph_pipe3;// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_ph_pipe4;// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_ph_pipe5;// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_ph_pipe6;// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_lp_ph_pipe7;// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fe_pipe0;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fe_pipe1;// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fe_pipe2;// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fe_pipe3;// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fe_pipe4;// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fe_pipe5;// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fe_pipe6;// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fe_pipe7;// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fs_pipe0;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fs_pipe1;// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fs_pipe2;// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fs_pipe3;// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fs_pipe4;// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fs_pipe5;// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fs_pipe6;// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_fs_pipe7;// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_le_pipe0;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_le_pipe1;// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_le_pipe2;// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_le_pipe3;// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_le_pipe4;// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_le_pipe5;// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_le_pipe6;// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_le_pipe7;// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_ls_pipe0;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_ls_pipe1;// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_ls_pipe2;// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_ls_pipe3;// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_ls_pipe4;// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_ls_pipe5;// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_ls_pipe6;// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_clear_resv_pkt_cnt_sp_ls_pipe7;// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [15:0]		reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input [15:0]		reg_dbg_pkt_num_nonzero_threshold;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input [9:0]		reg_dft_sync_tpram_config;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input [8:0]		reg_dft_tpram_config;	// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input			reg_last_byte_header_down_mux;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input			reg_resv_pkt_match_lp_dt_en_pipe0;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_resv_pkt_match_lp_dt_en_pipe1;// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_resv_pkt_match_lp_dt_en_pipe2;// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_resv_pkt_match_lp_dt_en_pipe3;// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_resv_pkt_match_lp_dt_en_pipe4;// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_resv_pkt_match_lp_dt_en_pipe5;// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_resv_pkt_match_lp_dt_en_pipe6;// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			reg_resv_pkt_match_lp_dt_en_pipe7;// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		reg_resv_pkt_match_lp_dt_pipe0;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		reg_resv_pkt_match_lp_dt_pipe1;// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		reg_resv_pkt_match_lp_dt_pipe2;// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		reg_resv_pkt_match_lp_dt_pipe3;// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		reg_resv_pkt_match_lp_dt_pipe4;// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		reg_resv_pkt_match_lp_dt_pipe5;// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		reg_resv_pkt_match_lp_dt_pipe6;// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [5:0]		reg_resv_pkt_match_lp_dt_pipe7;// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [7:0]		reg_sram_lcrc_err_oen;	// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input			reg_video_fifo_empty_depend_cnt_mux;// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input [7:0]		reg_video_pipe_en;	// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
input [16:0]		time_window0;		// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [16:0]		time_window1;		// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [16:0]		time_window2;		// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [16:0]		time_window3;		// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [16:0]		time_window4;		// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [16:0]		time_window5;		// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [16:0]		time_window6;		// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input [16:0]		time_window7;		// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			up_state_video_pipe0;	// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			up_state_video_pipe1;	// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			up_state_video_pipe2;	// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			up_state_video_pipe3;	// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			up_state_video_pipe4;	// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			up_state_video_pipe5;	// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			up_state_video_pipe6;	// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			up_state_video_pipe7;	// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			video_loss_en0;		// To u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			video_loss_en1;		// To u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			video_loss_en2;		// To u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			video_loss_en3;		// To u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			video_loss_en4;		// To u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			video_loss_en5;		// To u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			video_loss_en6;		// To u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
input			video_loss_en7;		// To u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
// End of automatics
input   [7:0]   pipe_fifo_full_clear;

/*AUTOOUTPUT*/
// Beginning of automatic outputs (from unused autoinst outputs)
output			ack0;			// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack1;			// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack2;			// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack3;			// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack4;			// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack5;			// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack6;			// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack7;			// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_pre0;		// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_pre1;		// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_pre2;		// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_pre3;		// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_pre4;		// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_pre5;		// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_pre6;		// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_pre7;		// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe0_aggregator0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe0_aggregator1;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe0_aggregator2;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe0_aggregator3;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe1_aggregator0;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe1_aggregator1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe1_aggregator2;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe1_aggregator3;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe2_aggregator0;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe2_aggregator1;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe2_aggregator2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe2_aggregator3;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe3_aggregator0;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe3_aggregator1;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe3_aggregator2;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe3_aggregator3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe4_aggregator0;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe4_aggregator1;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe4_aggregator2;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe4_aggregator3;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe5_aggregator0;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe5_aggregator1;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe5_aggregator2;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe5_aggregator3;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe6_aggregator0;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe6_aggregator1;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe6_aggregator2;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe6_aggregator3;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe7_aggregator0;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe7_aggregator1;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe7_aggregator2;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			ack_vld_pipe7_aggregator3;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe0_aggregator0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe0_aggregator1;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe0_aggregator2;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe0_aggregator3;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe1_aggregator0;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe1_aggregator1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe1_aggregator2;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe1_aggregator3;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe2_aggregator0;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe2_aggregator1;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe2_aggregator2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe2_aggregator3;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe3_aggregator0;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe3_aggregator1;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe3_aggregator2;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe3_aggregator3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe4_aggregator0;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe4_aggregator1;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe4_aggregator2;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe4_aggregator3;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe5_aggregator0;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe5_aggregator1;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe5_aggregator2;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe5_aggregator3;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe6_aggregator0;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe6_aggregator1;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe6_aggregator2;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe6_aggregator3;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe7_aggregator0;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe7_aggregator1;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe7_aggregator2;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			empty_vld_pipe7_aggregator3;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [2:0]		fifo_rd_ctrl_cs0;	// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [2:0]		fifo_rd_ctrl_cs1;	// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [2:0]		fifo_rd_ctrl_cs2;	// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [2:0]		fifo_rd_ctrl_cs3;	// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [2:0]		fifo_rd_ctrl_cs4;	// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [2:0]		fifo_rd_ctrl_cs5;	// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [2:0]		fifo_rd_ctrl_cs6;	// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [2:0]		fifo_rd_ctrl_cs7;	// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [15:0]		fs_cnt_pipe0;		// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [15:0]		fs_cnt_pipe1;		// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [15:0]		fs_cnt_pipe2;		// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [15:0]		fs_cnt_pipe3;		// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [15:0]		fs_cnt_pipe4;		// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [15:0]		fs_cnt_pipe5;		// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [15:0]		fs_cnt_pipe6;		// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [15:0]		fs_cnt_pipe7;		// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			fs_detect_pipe0;	// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			fs_detect_pipe1;	// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			fs_detect_pipe2;	// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			fs_detect_pipe3;	// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			fs_detect_pipe4;	// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			fs_detect_pipe5;	// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			fs_detect_pipe6;	// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			fs_detect_pipe7;	// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			lcrc_err0;		// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			lcrc_err1;		// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			lcrc_err2;		// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			lcrc_err3;		// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			lcrc_err4;		// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			lcrc_err5;		// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			lcrc_err6;		// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			lcrc_err7;		// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end0;		// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end1;		// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end2;		// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end3;		// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end4;		// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end5;		// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end6;		// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end7;		// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe0_aggregator0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe0_aggregator1;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe0_aggregator2;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe0_aggregator3;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe1_aggregator0;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe1_aggregator1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe1_aggregator2;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe1_aggregator3;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe2_aggregator0;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe2_aggregator1;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe2_aggregator2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe2_aggregator3;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe3_aggregator0;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe3_aggregator1;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe3_aggregator2;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe3_aggregator3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe4_aggregator0;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe4_aggregator1;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe4_aggregator2;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe4_aggregator3;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe5_aggregator0;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe5_aggregator1;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe5_aggregator2;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe5_aggregator3;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe6_aggregator0;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe6_aggregator1;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe6_aggregator2;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe6_aggregator3;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe7_aggregator0;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe7_aggregator1;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe7_aggregator2;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			line_end_vld_pipe7_aggregator3;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_async_fifo_pipe0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_async_fifo_pipe1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_async_fifo_pipe2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_async_fifo_pipe3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_async_fifo_pipe4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_async_fifo_pipe5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_async_fifo_pipe6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_async_fifo_pipe7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_sync_fifo_pipe0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_sync_fifo_pipe1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_sync_fifo_pipe2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_sync_fifo_pipe3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_sync_fifo_pipe4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_sync_fifo_pipe5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_sync_fifo_pipe6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_app_full_cnt_sync_fifo_pipe7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [7:0]		reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
output [7:0]		reg_rd_dbg_pkt_num_nonzero_threshold_err;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v, ...
output [31:0]		reg_rd_pipe0_dispatched_cnt_ready_for_sch;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_pipe1_dispatched_cnt_ready_for_sch;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_pipe2_dispatched_cnt_ready_for_sch;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_pipe3_dispatched_cnt_ready_for_sch;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_pipe4_dispatched_cnt_ready_for_sch;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_pipe5_dispatched_cnt_ready_for_sch;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_pipe6_dispatched_cnt_ready_for_sch;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_pipe7_dispatched_cnt_ready_for_sch;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_pf_pipe0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_pf_pipe1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_pf_pipe2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_pf_pipe3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_pf_pipe4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_pf_pipe5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_pf_pipe6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_pf_pipe7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_ph_pipe0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_ph_pipe1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_ph_pipe2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_ph_pipe3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_ph_pipe4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_ph_pipe5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_ph_pipe6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_lp_ph_pipe7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fe_pipe0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fe_pipe1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fe_pipe2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fe_pipe3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fe_pipe4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fe_pipe5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fe_pipe6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fe_pipe7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fs_pipe0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fs_pipe1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fs_pipe2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fs_pipe3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fs_pipe4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fs_pipe5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fs_pipe6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_fs_pipe7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_le_pipe0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_le_pipe1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_le_pipe2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_le_pipe3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_le_pipe4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_le_pipe5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_le_pipe6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_le_pipe7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_ls_pipe0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_ls_pipe1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_ls_pipe2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_ls_pipe3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_ls_pipe4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_ls_pipe5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_ls_pipe6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [31:0]		reg_rd_resv_pkt_cnt_sp_ls_pipe7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [(VIDEO_DATA_SIZE-1):0] video_data0;	// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [(VIDEO_DATA_SIZE-1):0] video_data1;	// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [(VIDEO_DATA_SIZE-1):0] video_data2;	// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [(VIDEO_DATA_SIZE-1):0] video_data3;	// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [(VIDEO_DATA_SIZE-1):0] video_data4;	// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [(VIDEO_DATA_SIZE-1):0] video_data5;	// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [(VIDEO_DATA_SIZE-1):0] video_data6;	// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [(VIDEO_DATA_SIZE-1):0] video_data7;	// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_double_err0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_double_err1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_double_err2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_double_err3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_double_err4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_double_err5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_double_err6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_double_err7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ecc_fault0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ecc_fault1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ecc_fault2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ecc_fault3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ecc_fault4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ecc_fault5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ecc_fault6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ecc_fault7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_empty0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_empty1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_empty2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_empty3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_empty4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_empty5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_empty6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_empty7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_full0;	// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_full1;	// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_full2;	// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_full3;	// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_full4;	// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_full5;	// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_full6;	// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_full7;	// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ovf_int0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ovf_int1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ovf_int2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ovf_int3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ovf_int4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ovf_int5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ovf_int6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_ovf_int7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_empty0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_empty1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_empty2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_empty3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_empty4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_empty5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_empty6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_empty7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_full0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_full1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_full2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_full3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_full4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_full5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_full6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_prog_full7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_single_err0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_single_err1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_single_err2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_single_err3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_single_err4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_single_err5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_single_err6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_single_err7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_udf_int0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_udf_int1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_udf_int2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_udf_int3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_udf_int4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_udf_int5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_udf_int6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_afifo_udf_int7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_double_err0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_double_err1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_double_err2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_double_err3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_double_err4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_double_err5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_double_err6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_double_err7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ecc_fault0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ecc_fault1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ecc_fault2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ecc_fault3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ecc_fault4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ecc_fault5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ecc_fault6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ecc_fault7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_empty0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_empty1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_empty2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_empty3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_empty4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_empty5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_empty6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_empty7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_full0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_full1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_full2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_full3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_full4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_full5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_full6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_full7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ovf_int0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ovf_int1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ovf_int2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ovf_int3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ovf_int4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ovf_int5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ovf_int6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_ovf_int7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_prog_full0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_prog_full1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_prog_full2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_prog_full3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_prog_full4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_prog_full5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_prog_full6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_prog_full7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_single_err0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_single_err1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_single_err2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_single_err3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_single_err4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_single_err5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_single_err6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_single_err7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_udf_int0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_udf_int1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_udf_int2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_udf_int3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_udf_int4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_udf_int5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_udf_int6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_fwft_fifo_udf_int7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_vld0;	// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_vld1;	// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_vld2;	// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_vld3;	// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_vld4;	// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_vld5;	// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_vld6;	// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_data_vld7;	// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_lock0;		// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_lock1;		// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_lock2;		// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_lock3;		// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_lock4;		// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_lock5;		// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_lock6;		// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_lock7;		// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_loss0;		// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_loss1;		// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_loss2;		// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_loss3;		// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_loss4;		// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_loss5;		// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_loss6;		// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_loss7;		// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [139:0]		video_pipe0_data_aggre_bypass;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe0_vld_aggre_bypass;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [139:0]		video_pipe1_data_aggre_bypass;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe1_vld_aggre_bypass;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [139:0]		video_pipe2_data_aggre_bypass;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe2_vld_aggre_bypass;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [139:0]		video_pipe3_data_aggre_bypass;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe3_vld_aggre_bypass;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [139:0]		video_pipe4_data_aggre_bypass;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe4_vld_aggre_bypass;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [139:0]		video_pipe5_data_aggre_bypass;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe5_vld_aggre_bypass;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [139:0]		video_pipe6_data_aggre_bypass;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe6_vld_aggre_bypass;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [139:0]		video_pipe7_data_aggre_bypass;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe7_vld_aggre_bypass;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [5:0]		video_pipe_date_type_for_concat_align0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [5:0]		video_pipe_date_type_for_concat_align1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [5:0]		video_pipe_date_type_for_concat_align2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [5:0]		video_pipe_date_type_for_concat_align3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [5:0]		video_pipe_date_type_for_concat_align4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [5:0]		video_pipe_date_type_for_concat_align5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [5:0]		video_pipe_date_type_for_concat_align6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output [5:0]		video_pipe_date_type_for_concat_align7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe_date_type_for_concat_align_vld0;// From u0_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe_date_type_for_concat_align_vld1;// From u1_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe_date_type_for_concat_align_vld2;// From u2_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe_date_type_for_concat_align_vld3;// From u3_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe_date_type_for_concat_align_vld4;// From u4_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe_date_type_for_concat_align_vld5;// From u5_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe_date_type_for_concat_align_vld6;// From u6_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
output			video_pipe_date_type_for_concat_align_vld7;// From u7_as6d_app_video_pipe_lane of as6d_app_video_pipe_lane.v
// End of automatics

output  [7:0]   reg_rd_pipe_fifo_full   ;


/*AUTOWIRE*/
// Beginning of automatic wires (for undeclared instantiated-module outputs)



//signal define pipe_fifo_full cnt
genvar          j                       ;
wire [7:0]      pipe_fifo_full_pre      ;
wire [7:0]      fifo_rdclk              ;
wire [7:0]      fifo_rdclk_rst_n        ;




 /*  as6d_app_video_pipe_lane  AUTO_TEMPLATE (
			.in_csi_data						(pipe@_csi_data[]),
			.in_bytes_en						(pipe@_bytes_en[]),
			.in_header_en						(pipe@_header_en),
			.in_data_en							(pipe@_data_en),
			.in_data_type						(pipe@_data_type[]),
			.in_virtual_channel					(pipe@_virtual_channel[]),
			.in_virtual_channel_x				(pipe@_virtual_channel_x[]),
			.in_word_count						(pipe@_word_count[]),
			.in_aggr_id							(pipe@_aggr_id[]),
			.in_pkt_crc					        (pipe@_pkt_crc[]),
			.in_pkt_crc_en				        (pipe@_pkt_crc_en[]),
			.up_state							(up_state_video_pipe@[]),
			.clk_1M								(clk_1M),
			.reg_dft_tpram_config				(reg_dft_tpram_config[]),
			.video_data_vld_aggregator\(.*\)	(pipe@_video_data_vld_aggregator\1[]),
			.reg_dft_sync_tpram_config			(reg_dft_sync_tpram_config[]),
			.empty_vld_aggregator0				(empty_vld_pipe@_aggregator0),
			.empty_vld_aggregator1				(empty_vld_pipe@_aggregator1),
			.empty_vld_aggregator2				(empty_vld_pipe@_aggregator2),
			.empty_vld_aggregator3				(empty_vld_pipe@_aggregator3),
			.ack_vld_aggregator0				(ack_vld_pipe@_aggregator0),
			.ack_vld_aggregator1				(ack_vld_pipe@_aggregator1),
			.ack_vld_aggregator2				(ack_vld_pipe@_aggregator2),
			.ack_vld_aggregator3				(ack_vld_pipe@_aggregator3),
			.line_end_vld_aggregator0			(line_end_vld_pipe@_aggregator0),
			.line_end_vld_aggregator1			(line_end_vld_pipe@_aggregator1),
			.line_end_vld_aggregator2			(line_end_vld_pipe@_aggregator2),
			.line_end_vld_aggregator3			(line_end_vld_pipe@_aggregator3),
			.app_aggregation_bypass             (app_aggregation_bypass),
			.video_pipe_data_aggre_bypass       (video_pipe@_data_aggre_bypass[139:0]),
			.video_pipe_vld_aggre_bypass        (video_pipe@_vld_aggre_bypass),
			.reg_rd_resv_\(.*\)                 (reg_rd_resv_\1_pipe@[]), 
			.reg_resv_\(.*\)                 (reg_resv_\1_pipe@[]), 
            .reg_clear_resv_\(.*\)              (reg_clear_resv_\1_pipe@[]),
			.reg_video_fifo_empty_depend_cnt_mux(reg_video_fifo_empty_depend_cnt_mux),
			.reg_last_byte_header_down_mux(reg_last_byte_header_down_mux),
			.reg_rd_resv_\(.*\)                 (reg_rd_resv_\1_pipe@[]), 
            .reg_clear_resv_\(.*\)              (reg_clear_resv_\1_pipe@[]),
			.reg_rd_app_\(.*\)                  (reg_rd_app_\1_pipe@[]), 
			.reg_clear_app_\(.*\)               (reg_clear_app_\1_pipe@[]), 
			.reg_rd_dispatched_cnt_ready_for_sch(reg_rd_pipe@_dispatched_cnt_ready_for_sch[]), 
			.reg_app_pkt_crc_gen_dis(reg_app_pkt_crc_gen_dis),
			.reg_sram_lcrc_err_oen(reg_sram_lcrc_err_oen[@]),
			.reg_video_pipe_en(reg_video_pipe_en[@]),
			.reg_app_ecc_addr_protect_en(reg_app_ecc_addr_protect_en),
			.reg_app_ecc_bypass(reg_app_ecc_bypass),
			.reg_app_ecc_fault_detc_en(reg_app_ecc_fault_detc_en),
			.reg_app_wr_idi_data_continue(reg_app_wr_idi_data_continue),
            .reg_rd_dbg_pkt_num_nonzero_threshold_err(reg_rd_dbg_pkt_num_nonzero_threshold_err[@]),
            .reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err(reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err[@]),
            .reg_dbg_pkt_num_nonzero_threshold(reg_dbg_pkt_num_nonzero_threshold[]),
            .reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold(reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold[]),
            .\(.*\)   (\1@[]),

 ) */
as6d_app_video_pipe_lane    u0_as6d_app_video_pipe_lane(/*AUTOINST*/
							// Outputs
							.ack_pre	(ack_pre0),	 // Templated
							.video_data_afifo_ecc_fault(video_data_afifo_ecc_fault0), // Templated
							.video_data_fwft_fifo_ecc_fault(video_data_fwft_fifo_ecc_fault0), // Templated
							.video_data_afifo_single_err(video_data_afifo_single_err0), // Templated
							.video_data_afifo_double_err(video_data_afifo_double_err0), // Templated
							.video_data_afifo_ovf_int(video_data_afifo_ovf_int0), // Templated
							.video_data_afifo_udf_int(video_data_afifo_udf_int0), // Templated
							.video_data_afifo_prog_full(video_data_afifo_prog_full0), // Templated
							.video_data_afifo_empty(video_data_afifo_empty0), // Templated
							.video_data_afifo_full(video_data_afifo_full0), // Templated
							.video_data_afifo_prog_empty(video_data_afifo_prog_empty0), // Templated
							.video_data_fwft_fifo_single_err(video_data_fwft_fifo_single_err0), // Templated
							.video_data_fwft_fifo_double_err(video_data_fwft_fifo_double_err0), // Templated
							.video_data_fwft_fifo_ovf_int(video_data_fwft_fifo_ovf_int0), // Templated
							.video_data_fwft_fifo_udf_int(video_data_fwft_fifo_udf_int0), // Templated
							.video_data_fwft_fifo_prog_full(video_data_fwft_fifo_prog_full0), // Templated
							.video_data_fwft_fifo_empty(video_data_fwft_fifo_empty0), // Templated
							.video_data_fwft_fifo_full(video_data_fwft_fifo_full0), // Templated
							.video_data_vld	(video_data_vld0), // Templated
							.video_data	(video_data0[(VIDEO_DATA_SIZE-1):0]), // Templated
							.ack		(ack0),		 // Templated
							.line_end	(line_end0),	 // Templated
							.video_loss	(video_loss0),	 // Templated
							.video_lock	(video_lock0),	 // Templated
							.fifo_rd_ctrl_cs(fifo_rd_ctrl_cs0[2:0]), // Templated
							.fs_detect_pipe	(fs_detect_pipe0), // Templated
							.fs_cnt_pipe	(fs_cnt_pipe0[15:0]), // Templated
							.empty_vld_aggregator0(empty_vld_pipe0_aggregator0), // Templated
							.empty_vld_aggregator1(empty_vld_pipe0_aggregator1), // Templated
							.empty_vld_aggregator2(empty_vld_pipe0_aggregator2), // Templated
							.empty_vld_aggregator3(empty_vld_pipe0_aggregator3), // Templated
							.ack_vld_aggregator0(ack_vld_pipe0_aggregator0), // Templated
							.ack_vld_aggregator1(ack_vld_pipe0_aggregator1), // Templated
							.ack_vld_aggregator2(ack_vld_pipe0_aggregator2), // Templated
							.ack_vld_aggregator3(ack_vld_pipe0_aggregator3), // Templated
							.line_end_vld_aggregator0(line_end_vld_pipe0_aggregator0), // Templated
							.line_end_vld_aggregator1(line_end_vld_pipe0_aggregator1), // Templated
							.line_end_vld_aggregator2(line_end_vld_pipe0_aggregator2), // Templated
							.line_end_vld_aggregator3(line_end_vld_pipe0_aggregator3), // Templated
							.video_pipe_data_aggre_bypass(video_pipe0_data_aggre_bypass[139:0]), // Templated
							.video_pipe_vld_aggre_bypass(video_pipe0_vld_aggre_bypass), // Templated
							.reg_rd_resv_pkt_cnt_lp_pf(reg_rd_resv_pkt_cnt_lp_pf_pipe0[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_lp_ph(reg_rd_resv_pkt_cnt_lp_ph_pipe0[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_le(reg_rd_resv_pkt_cnt_sp_le_pipe0[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_ls(reg_rd_resv_pkt_cnt_sp_ls_pipe0[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fe(reg_rd_resv_pkt_cnt_sp_fe_pipe0[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fs(reg_rd_resv_pkt_cnt_sp_fs_pipe0[31:0]), // Templated
							.reg_rd_app_full_cnt_sync_fifo(reg_rd_app_full_cnt_sync_fifo_pipe0[31:0]), // Templated
							.reg_rd_app_full_cnt_async_fifo(reg_rd_app_full_cnt_async_fifo_pipe0[31:0]), // Templated
							.reg_rd_dispatched_cnt_ready_for_sch(reg_rd_pipe0_dispatched_cnt_ready_for_sch[31:0]), // Templated
							.lcrc_err	(lcrc_err0),	 // Templated
							.reg_rd_dbg_pkt_num_nonzero_threshold_err(reg_rd_dbg_pkt_num_nonzero_threshold_err[0]), // Templated
							.reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err(reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err[0]), // Templated
							.video_pipe_date_type_for_concat_align(video_pipe_date_type_for_concat_align0[5:0]), // Templated
							.video_pipe_date_type_for_concat_align_vld(video_pipe_date_type_for_concat_align_vld0), // Templated
							// Inputs
							.reg_app_ecc_addr_protect_en(reg_app_ecc_addr_protect_en), // Templated
							.reg_app_ecc_bypass(reg_app_ecc_bypass), // Templated
							.reg_app_ecc_fault_detc_en(reg_app_ecc_fault_detc_en), // Templated
							.reg_app_pkt_crc_gen_dis(reg_app_pkt_crc_gen_dis), // Templated
							.reg_resv_pkt_match_lp_dt(reg_resv_pkt_match_lp_dt_pipe0[5:0]), // Templated
							.reg_resv_pkt_match_lp_dt_en(reg_resv_pkt_match_lp_dt_en_pipe0), // Templated
							.reg_sram_lcrc_err_oen(reg_sram_lcrc_err_oen[0]), // Templated
							.reg_video_fifo_empty_depend_cnt_mux(reg_video_fifo_empty_depend_cnt_mux), // Templated
							.clk_1M		(clk_1M),	 // Templated
							.fifo_wrclk	(fifo_wrclk0),	 // Templated
							.fifo_wrclk_rst_n(fifo_wrclk_rst_n0), // Templated
							.fifo_rdclk	(fifo_rdclk0),	 // Templated
							.fifo_rdclk_rst_n(fifo_rdclk_rst_n0), // Templated
							.in_csi_data	(pipe0_csi_data[(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0]), // Templated
							.in_bytes_en	(pipe0_bytes_en[(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0]), // Templated
							.in_header_en	(pipe0_header_en), // Templated
							.in_data_en	(pipe0_data_en), // Templated
							.in_data_type	(pipe0_data_type[5:0]), // Templated
							.in_virtual_channel(pipe0_virtual_channel[1:0]), // Templated
							.in_virtual_channel_x(pipe0_virtual_channel_x[(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0]), // Templated
							.in_word_count	(pipe0_word_count[15:0]), // Templated
							.in_aggr_id	(pipe0_aggr_id[3:0]), // Templated
							.in_pkt_crc	(pipe0_pkt_crc[31:0]), // Templated
							.in_pkt_crc_en	(pipe0_pkt_crc_en), // Templated
							.up_state	(up_state_video_pipe0), // Templated
							.line_delay_en	(line_delay_en0), // Templated
							.video_loss_en	(video_loss_en0), // Templated
							.time_window	(time_window0[16:0]), // Templated
							.reg_dft_tpram_config(reg_dft_tpram_config[8:0]), // Templated
							.reg_dft_sync_tpram_config(reg_dft_sync_tpram_config[9:0]), // Templated
							.app_aggregation_bypass(app_aggregation_bypass), // Templated
							.reg_video_pipe_en(reg_video_pipe_en[0]), // Templated
							.reg_last_byte_header_down_mux(reg_last_byte_header_down_mux), // Templated
							.reg_clear_resv_pkt_cnt_lp_pf(reg_clear_resv_pkt_cnt_lp_pf_pipe0), // Templated
							.reg_clear_resv_pkt_cnt_lp_ph(reg_clear_resv_pkt_cnt_lp_ph_pipe0), // Templated
							.reg_clear_resv_pkt_cnt_sp_le(reg_clear_resv_pkt_cnt_sp_le_pipe0), // Templated
							.reg_clear_resv_pkt_cnt_sp_ls(reg_clear_resv_pkt_cnt_sp_ls_pipe0), // Templated
							.reg_clear_resv_pkt_cnt_sp_fe(reg_clear_resv_pkt_cnt_sp_fe_pipe0), // Templated
							.reg_clear_resv_pkt_cnt_sp_fs(reg_clear_resv_pkt_cnt_sp_fs_pipe0), // Templated
							.reg_clear_app_full_cnt_async_fifo(reg_clear_app_full_cnt_async_fifo_pipe0), // Templated
							.reg_clear_app_full_cnt_sync_fifo(reg_clear_app_full_cnt_sync_fifo_pipe0), // Templated
							.reg_app_wr_idi_data_continue(reg_app_wr_idi_data_continue), // Templated
							.reg_dbg_pkt_num_nonzero_threshold(reg_dbg_pkt_num_nonzero_threshold[15:0]), // Templated
							.reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold(reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold[15:0])); // Templated


as6d_app_video_pipe_lane    u1_as6d_app_video_pipe_lane(/*AUTOINST*/
							// Outputs
							.ack_pre	(ack_pre1),	 // Templated
							.video_data_afifo_ecc_fault(video_data_afifo_ecc_fault1), // Templated
							.video_data_fwft_fifo_ecc_fault(video_data_fwft_fifo_ecc_fault1), // Templated
							.video_data_afifo_single_err(video_data_afifo_single_err1), // Templated
							.video_data_afifo_double_err(video_data_afifo_double_err1), // Templated
							.video_data_afifo_ovf_int(video_data_afifo_ovf_int1), // Templated
							.video_data_afifo_udf_int(video_data_afifo_udf_int1), // Templated
							.video_data_afifo_prog_full(video_data_afifo_prog_full1), // Templated
							.video_data_afifo_empty(video_data_afifo_empty1), // Templated
							.video_data_afifo_full(video_data_afifo_full1), // Templated
							.video_data_afifo_prog_empty(video_data_afifo_prog_empty1), // Templated
							.video_data_fwft_fifo_single_err(video_data_fwft_fifo_single_err1), // Templated
							.video_data_fwft_fifo_double_err(video_data_fwft_fifo_double_err1), // Templated
							.video_data_fwft_fifo_ovf_int(video_data_fwft_fifo_ovf_int1), // Templated
							.video_data_fwft_fifo_udf_int(video_data_fwft_fifo_udf_int1), // Templated
							.video_data_fwft_fifo_prog_full(video_data_fwft_fifo_prog_full1), // Templated
							.video_data_fwft_fifo_empty(video_data_fwft_fifo_empty1), // Templated
							.video_data_fwft_fifo_full(video_data_fwft_fifo_full1), // Templated
							.video_data_vld	(video_data_vld1), // Templated
							.video_data	(video_data1[(VIDEO_DATA_SIZE-1):0]), // Templated
							.ack		(ack1),		 // Templated
							.line_end	(line_end1),	 // Templated
							.video_loss	(video_loss1),	 // Templated
							.video_lock	(video_lock1),	 // Templated
							.fifo_rd_ctrl_cs(fifo_rd_ctrl_cs1[2:0]), // Templated
							.fs_detect_pipe	(fs_detect_pipe1), // Templated
							.fs_cnt_pipe	(fs_cnt_pipe1[15:0]), // Templated
							.empty_vld_aggregator0(empty_vld_pipe1_aggregator0), // Templated
							.empty_vld_aggregator1(empty_vld_pipe1_aggregator1), // Templated
							.empty_vld_aggregator2(empty_vld_pipe1_aggregator2), // Templated
							.empty_vld_aggregator3(empty_vld_pipe1_aggregator3), // Templated
							.ack_vld_aggregator0(ack_vld_pipe1_aggregator0), // Templated
							.ack_vld_aggregator1(ack_vld_pipe1_aggregator1), // Templated
							.ack_vld_aggregator2(ack_vld_pipe1_aggregator2), // Templated
							.ack_vld_aggregator3(ack_vld_pipe1_aggregator3), // Templated
							.line_end_vld_aggregator0(line_end_vld_pipe1_aggregator0), // Templated
							.line_end_vld_aggregator1(line_end_vld_pipe1_aggregator1), // Templated
							.line_end_vld_aggregator2(line_end_vld_pipe1_aggregator2), // Templated
							.line_end_vld_aggregator3(line_end_vld_pipe1_aggregator3), // Templated
							.video_pipe_data_aggre_bypass(video_pipe1_data_aggre_bypass[139:0]), // Templated
							.video_pipe_vld_aggre_bypass(video_pipe1_vld_aggre_bypass), // Templated
							.reg_rd_resv_pkt_cnt_lp_pf(reg_rd_resv_pkt_cnt_lp_pf_pipe1[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_lp_ph(reg_rd_resv_pkt_cnt_lp_ph_pipe1[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_le(reg_rd_resv_pkt_cnt_sp_le_pipe1[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_ls(reg_rd_resv_pkt_cnt_sp_ls_pipe1[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fe(reg_rd_resv_pkt_cnt_sp_fe_pipe1[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fs(reg_rd_resv_pkt_cnt_sp_fs_pipe1[31:0]), // Templated
							.reg_rd_app_full_cnt_sync_fifo(reg_rd_app_full_cnt_sync_fifo_pipe1[31:0]), // Templated
							.reg_rd_app_full_cnt_async_fifo(reg_rd_app_full_cnt_async_fifo_pipe1[31:0]), // Templated
							.reg_rd_dispatched_cnt_ready_for_sch(reg_rd_pipe1_dispatched_cnt_ready_for_sch[31:0]), // Templated
							.lcrc_err	(lcrc_err1),	 // Templated
							.reg_rd_dbg_pkt_num_nonzero_threshold_err(reg_rd_dbg_pkt_num_nonzero_threshold_err[1]), // Templated
							.reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err(reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err[1]), // Templated
							.video_pipe_date_type_for_concat_align(video_pipe_date_type_for_concat_align1[5:0]), // Templated
							.video_pipe_date_type_for_concat_align_vld(video_pipe_date_type_for_concat_align_vld1), // Templated
							// Inputs
							.reg_app_ecc_addr_protect_en(reg_app_ecc_addr_protect_en), // Templated
							.reg_app_ecc_bypass(reg_app_ecc_bypass), // Templated
							.reg_app_ecc_fault_detc_en(reg_app_ecc_fault_detc_en), // Templated
							.reg_app_pkt_crc_gen_dis(reg_app_pkt_crc_gen_dis), // Templated
							.reg_resv_pkt_match_lp_dt(reg_resv_pkt_match_lp_dt_pipe1[5:0]), // Templated
							.reg_resv_pkt_match_lp_dt_en(reg_resv_pkt_match_lp_dt_en_pipe1), // Templated
							.reg_sram_lcrc_err_oen(reg_sram_lcrc_err_oen[1]), // Templated
							.reg_video_fifo_empty_depend_cnt_mux(reg_video_fifo_empty_depend_cnt_mux), // Templated
							.clk_1M		(clk_1M),	 // Templated
							.fifo_wrclk	(fifo_wrclk1),	 // Templated
							.fifo_wrclk_rst_n(fifo_wrclk_rst_n1), // Templated
							.fifo_rdclk	(fifo_rdclk1),	 // Templated
							.fifo_rdclk_rst_n(fifo_rdclk_rst_n1), // Templated
							.in_csi_data	(pipe1_csi_data[(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0]), // Templated
							.in_bytes_en	(pipe1_bytes_en[(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0]), // Templated
							.in_header_en	(pipe1_header_en), // Templated
							.in_data_en	(pipe1_data_en), // Templated
							.in_data_type	(pipe1_data_type[5:0]), // Templated
							.in_virtual_channel(pipe1_virtual_channel[1:0]), // Templated
							.in_virtual_channel_x(pipe1_virtual_channel_x[(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0]), // Templated
							.in_word_count	(pipe1_word_count[15:0]), // Templated
							.in_aggr_id	(pipe1_aggr_id[3:0]), // Templated
							.in_pkt_crc	(pipe1_pkt_crc[31:0]), // Templated
							.in_pkt_crc_en	(pipe1_pkt_crc_en), // Templated
							.up_state	(up_state_video_pipe1), // Templated
							.line_delay_en	(line_delay_en1), // Templated
							.video_loss_en	(video_loss_en1), // Templated
							.time_window	(time_window1[16:0]), // Templated
							.reg_dft_tpram_config(reg_dft_tpram_config[8:0]), // Templated
							.reg_dft_sync_tpram_config(reg_dft_sync_tpram_config[9:0]), // Templated
							.app_aggregation_bypass(app_aggregation_bypass), // Templated
							.reg_video_pipe_en(reg_video_pipe_en[1]), // Templated
							.reg_last_byte_header_down_mux(reg_last_byte_header_down_mux), // Templated
							.reg_clear_resv_pkt_cnt_lp_pf(reg_clear_resv_pkt_cnt_lp_pf_pipe1), // Templated
							.reg_clear_resv_pkt_cnt_lp_ph(reg_clear_resv_pkt_cnt_lp_ph_pipe1), // Templated
							.reg_clear_resv_pkt_cnt_sp_le(reg_clear_resv_pkt_cnt_sp_le_pipe1), // Templated
							.reg_clear_resv_pkt_cnt_sp_ls(reg_clear_resv_pkt_cnt_sp_ls_pipe1), // Templated
							.reg_clear_resv_pkt_cnt_sp_fe(reg_clear_resv_pkt_cnt_sp_fe_pipe1), // Templated
							.reg_clear_resv_pkt_cnt_sp_fs(reg_clear_resv_pkt_cnt_sp_fs_pipe1), // Templated
							.reg_clear_app_full_cnt_async_fifo(reg_clear_app_full_cnt_async_fifo_pipe1), // Templated
							.reg_clear_app_full_cnt_sync_fifo(reg_clear_app_full_cnt_sync_fifo_pipe1), // Templated
							.reg_app_wr_idi_data_continue(reg_app_wr_idi_data_continue), // Templated
							.reg_dbg_pkt_num_nonzero_threshold(reg_dbg_pkt_num_nonzero_threshold[15:0]), // Templated
							.reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold(reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold[15:0])); // Templated
as6d_app_video_pipe_lane    u2_as6d_app_video_pipe_lane(/*AUTOINST*/
							// Outputs
							.ack_pre	(ack_pre2),	 // Templated
							.video_data_afifo_ecc_fault(video_data_afifo_ecc_fault2), // Templated
							.video_data_fwft_fifo_ecc_fault(video_data_fwft_fifo_ecc_fault2), // Templated
							.video_data_afifo_single_err(video_data_afifo_single_err2), // Templated
							.video_data_afifo_double_err(video_data_afifo_double_err2), // Templated
							.video_data_afifo_ovf_int(video_data_afifo_ovf_int2), // Templated
							.video_data_afifo_udf_int(video_data_afifo_udf_int2), // Templated
							.video_data_afifo_prog_full(video_data_afifo_prog_full2), // Templated
							.video_data_afifo_empty(video_data_afifo_empty2), // Templated
							.video_data_afifo_full(video_data_afifo_full2), // Templated
							.video_data_afifo_prog_empty(video_data_afifo_prog_empty2), // Templated
							.video_data_fwft_fifo_single_err(video_data_fwft_fifo_single_err2), // Templated
							.video_data_fwft_fifo_double_err(video_data_fwft_fifo_double_err2), // Templated
							.video_data_fwft_fifo_ovf_int(video_data_fwft_fifo_ovf_int2), // Templated
							.video_data_fwft_fifo_udf_int(video_data_fwft_fifo_udf_int2), // Templated
							.video_data_fwft_fifo_prog_full(video_data_fwft_fifo_prog_full2), // Templated
							.video_data_fwft_fifo_empty(video_data_fwft_fifo_empty2), // Templated
							.video_data_fwft_fifo_full(video_data_fwft_fifo_full2), // Templated
							.video_data_vld	(video_data_vld2), // Templated
							.video_data	(video_data2[(VIDEO_DATA_SIZE-1):0]), // Templated
							.ack		(ack2),		 // Templated
							.line_end	(line_end2),	 // Templated
							.video_loss	(video_loss2),	 // Templated
							.video_lock	(video_lock2),	 // Templated
							.fifo_rd_ctrl_cs(fifo_rd_ctrl_cs2[2:0]), // Templated
							.fs_detect_pipe	(fs_detect_pipe2), // Templated
							.fs_cnt_pipe	(fs_cnt_pipe2[15:0]), // Templated
							.empty_vld_aggregator0(empty_vld_pipe2_aggregator0), // Templated
							.empty_vld_aggregator1(empty_vld_pipe2_aggregator1), // Templated
							.empty_vld_aggregator2(empty_vld_pipe2_aggregator2), // Templated
							.empty_vld_aggregator3(empty_vld_pipe2_aggregator3), // Templated
							.ack_vld_aggregator0(ack_vld_pipe2_aggregator0), // Templated
							.ack_vld_aggregator1(ack_vld_pipe2_aggregator1), // Templated
							.ack_vld_aggregator2(ack_vld_pipe2_aggregator2), // Templated
							.ack_vld_aggregator3(ack_vld_pipe2_aggregator3), // Templated
							.line_end_vld_aggregator0(line_end_vld_pipe2_aggregator0), // Templated
							.line_end_vld_aggregator1(line_end_vld_pipe2_aggregator1), // Templated
							.line_end_vld_aggregator2(line_end_vld_pipe2_aggregator2), // Templated
							.line_end_vld_aggregator3(line_end_vld_pipe2_aggregator3), // Templated
							.video_pipe_data_aggre_bypass(video_pipe2_data_aggre_bypass[139:0]), // Templated
							.video_pipe_vld_aggre_bypass(video_pipe2_vld_aggre_bypass), // Templated
							.reg_rd_resv_pkt_cnt_lp_pf(reg_rd_resv_pkt_cnt_lp_pf_pipe2[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_lp_ph(reg_rd_resv_pkt_cnt_lp_ph_pipe2[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_le(reg_rd_resv_pkt_cnt_sp_le_pipe2[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_ls(reg_rd_resv_pkt_cnt_sp_ls_pipe2[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fe(reg_rd_resv_pkt_cnt_sp_fe_pipe2[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fs(reg_rd_resv_pkt_cnt_sp_fs_pipe2[31:0]), // Templated
							.reg_rd_app_full_cnt_sync_fifo(reg_rd_app_full_cnt_sync_fifo_pipe2[31:0]), // Templated
							.reg_rd_app_full_cnt_async_fifo(reg_rd_app_full_cnt_async_fifo_pipe2[31:0]), // Templated
							.reg_rd_dispatched_cnt_ready_for_sch(reg_rd_pipe2_dispatched_cnt_ready_for_sch[31:0]), // Templated
							.lcrc_err	(lcrc_err2),	 // Templated
							.reg_rd_dbg_pkt_num_nonzero_threshold_err(reg_rd_dbg_pkt_num_nonzero_threshold_err[2]), // Templated
							.reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err(reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err[2]), // Templated
							.video_pipe_date_type_for_concat_align(video_pipe_date_type_for_concat_align2[5:0]), // Templated
							.video_pipe_date_type_for_concat_align_vld(video_pipe_date_type_for_concat_align_vld2), // Templated
							// Inputs
							.reg_app_ecc_addr_protect_en(reg_app_ecc_addr_protect_en), // Templated
							.reg_app_ecc_bypass(reg_app_ecc_bypass), // Templated
							.reg_app_ecc_fault_detc_en(reg_app_ecc_fault_detc_en), // Templated
							.reg_app_pkt_crc_gen_dis(reg_app_pkt_crc_gen_dis), // Templated
							.reg_resv_pkt_match_lp_dt(reg_resv_pkt_match_lp_dt_pipe2[5:0]), // Templated
							.reg_resv_pkt_match_lp_dt_en(reg_resv_pkt_match_lp_dt_en_pipe2), // Templated
							.reg_sram_lcrc_err_oen(reg_sram_lcrc_err_oen[2]), // Templated
							.reg_video_fifo_empty_depend_cnt_mux(reg_video_fifo_empty_depend_cnt_mux), // Templated
							.clk_1M		(clk_1M),	 // Templated
							.fifo_wrclk	(fifo_wrclk2),	 // Templated
							.fifo_wrclk_rst_n(fifo_wrclk_rst_n2), // Templated
							.fifo_rdclk	(fifo_rdclk2),	 // Templated
							.fifo_rdclk_rst_n(fifo_rdclk_rst_n2), // Templated
							.in_csi_data	(pipe2_csi_data[(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0]), // Templated
							.in_bytes_en	(pipe2_bytes_en[(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0]), // Templated
							.in_header_en	(pipe2_header_en), // Templated
							.in_data_en	(pipe2_data_en), // Templated
							.in_data_type	(pipe2_data_type[5:0]), // Templated
							.in_virtual_channel(pipe2_virtual_channel[1:0]), // Templated
							.in_virtual_channel_x(pipe2_virtual_channel_x[(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0]), // Templated
							.in_word_count	(pipe2_word_count[15:0]), // Templated
							.in_aggr_id	(pipe2_aggr_id[3:0]), // Templated
							.in_pkt_crc	(pipe2_pkt_crc[31:0]), // Templated
							.in_pkt_crc_en	(pipe2_pkt_crc_en), // Templated
							.up_state	(up_state_video_pipe2), // Templated
							.line_delay_en	(line_delay_en2), // Templated
							.video_loss_en	(video_loss_en2), // Templated
							.time_window	(time_window2[16:0]), // Templated
							.reg_dft_tpram_config(reg_dft_tpram_config[8:0]), // Templated
							.reg_dft_sync_tpram_config(reg_dft_sync_tpram_config[9:0]), // Templated
							.app_aggregation_bypass(app_aggregation_bypass), // Templated
							.reg_video_pipe_en(reg_video_pipe_en[2]), // Templated
							.reg_last_byte_header_down_mux(reg_last_byte_header_down_mux), // Templated
							.reg_clear_resv_pkt_cnt_lp_pf(reg_clear_resv_pkt_cnt_lp_pf_pipe2), // Templated
							.reg_clear_resv_pkt_cnt_lp_ph(reg_clear_resv_pkt_cnt_lp_ph_pipe2), // Templated
							.reg_clear_resv_pkt_cnt_sp_le(reg_clear_resv_pkt_cnt_sp_le_pipe2), // Templated
							.reg_clear_resv_pkt_cnt_sp_ls(reg_clear_resv_pkt_cnt_sp_ls_pipe2), // Templated
							.reg_clear_resv_pkt_cnt_sp_fe(reg_clear_resv_pkt_cnt_sp_fe_pipe2), // Templated
							.reg_clear_resv_pkt_cnt_sp_fs(reg_clear_resv_pkt_cnt_sp_fs_pipe2), // Templated
							.reg_clear_app_full_cnt_async_fifo(reg_clear_app_full_cnt_async_fifo_pipe2), // Templated
							.reg_clear_app_full_cnt_sync_fifo(reg_clear_app_full_cnt_sync_fifo_pipe2), // Templated
							.reg_app_wr_idi_data_continue(reg_app_wr_idi_data_continue), // Templated
							.reg_dbg_pkt_num_nonzero_threshold(reg_dbg_pkt_num_nonzero_threshold[15:0]), // Templated
							.reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold(reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold[15:0])); // Templated
as6d_app_video_pipe_lane    u3_as6d_app_video_pipe_lane(/*AUTOINST*/
							// Outputs
							.ack_pre	(ack_pre3),	 // Templated
							.video_data_afifo_ecc_fault(video_data_afifo_ecc_fault3), // Templated
							.video_data_fwft_fifo_ecc_fault(video_data_fwft_fifo_ecc_fault3), // Templated
							.video_data_afifo_single_err(video_data_afifo_single_err3), // Templated
							.video_data_afifo_double_err(video_data_afifo_double_err3), // Templated
							.video_data_afifo_ovf_int(video_data_afifo_ovf_int3), // Templated
							.video_data_afifo_udf_int(video_data_afifo_udf_int3), // Templated
							.video_data_afifo_prog_full(video_data_afifo_prog_full3), // Templated
							.video_data_afifo_empty(video_data_afifo_empty3), // Templated
							.video_data_afifo_full(video_data_afifo_full3), // Templated
							.video_data_afifo_prog_empty(video_data_afifo_prog_empty3), // Templated
							.video_data_fwft_fifo_single_err(video_data_fwft_fifo_single_err3), // Templated
							.video_data_fwft_fifo_double_err(video_data_fwft_fifo_double_err3), // Templated
							.video_data_fwft_fifo_ovf_int(video_data_fwft_fifo_ovf_int3), // Templated
							.video_data_fwft_fifo_udf_int(video_data_fwft_fifo_udf_int3), // Templated
							.video_data_fwft_fifo_prog_full(video_data_fwft_fifo_prog_full3), // Templated
							.video_data_fwft_fifo_empty(video_data_fwft_fifo_empty3), // Templated
							.video_data_fwft_fifo_full(video_data_fwft_fifo_full3), // Templated
							.video_data_vld	(video_data_vld3), // Templated
							.video_data	(video_data3[(VIDEO_DATA_SIZE-1):0]), // Templated
							.ack		(ack3),		 // Templated
							.line_end	(line_end3),	 // Templated
							.video_loss	(video_loss3),	 // Templated
							.video_lock	(video_lock3),	 // Templated
							.fifo_rd_ctrl_cs(fifo_rd_ctrl_cs3[2:0]), // Templated
							.fs_detect_pipe	(fs_detect_pipe3), // Templated
							.fs_cnt_pipe	(fs_cnt_pipe3[15:0]), // Templated
							.empty_vld_aggregator0(empty_vld_pipe3_aggregator0), // Templated
							.empty_vld_aggregator1(empty_vld_pipe3_aggregator1), // Templated
							.empty_vld_aggregator2(empty_vld_pipe3_aggregator2), // Templated
							.empty_vld_aggregator3(empty_vld_pipe3_aggregator3), // Templated
							.ack_vld_aggregator0(ack_vld_pipe3_aggregator0), // Templated
							.ack_vld_aggregator1(ack_vld_pipe3_aggregator1), // Templated
							.ack_vld_aggregator2(ack_vld_pipe3_aggregator2), // Templated
							.ack_vld_aggregator3(ack_vld_pipe3_aggregator3), // Templated
							.line_end_vld_aggregator0(line_end_vld_pipe3_aggregator0), // Templated
							.line_end_vld_aggregator1(line_end_vld_pipe3_aggregator1), // Templated
							.line_end_vld_aggregator2(line_end_vld_pipe3_aggregator2), // Templated
							.line_end_vld_aggregator3(line_end_vld_pipe3_aggregator3), // Templated
							.video_pipe_data_aggre_bypass(video_pipe3_data_aggre_bypass[139:0]), // Templated
							.video_pipe_vld_aggre_bypass(video_pipe3_vld_aggre_bypass), // Templated
							.reg_rd_resv_pkt_cnt_lp_pf(reg_rd_resv_pkt_cnt_lp_pf_pipe3[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_lp_ph(reg_rd_resv_pkt_cnt_lp_ph_pipe3[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_le(reg_rd_resv_pkt_cnt_sp_le_pipe3[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_ls(reg_rd_resv_pkt_cnt_sp_ls_pipe3[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fe(reg_rd_resv_pkt_cnt_sp_fe_pipe3[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fs(reg_rd_resv_pkt_cnt_sp_fs_pipe3[31:0]), // Templated
							.reg_rd_app_full_cnt_sync_fifo(reg_rd_app_full_cnt_sync_fifo_pipe3[31:0]), // Templated
							.reg_rd_app_full_cnt_async_fifo(reg_rd_app_full_cnt_async_fifo_pipe3[31:0]), // Templated
							.reg_rd_dispatched_cnt_ready_for_sch(reg_rd_pipe3_dispatched_cnt_ready_for_sch[31:0]), // Templated
							.lcrc_err	(lcrc_err3),	 // Templated
							.reg_rd_dbg_pkt_num_nonzero_threshold_err(reg_rd_dbg_pkt_num_nonzero_threshold_err[3]), // Templated
							.reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err(reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err[3]), // Templated
							.video_pipe_date_type_for_concat_align(video_pipe_date_type_for_concat_align3[5:0]), // Templated
							.video_pipe_date_type_for_concat_align_vld(video_pipe_date_type_for_concat_align_vld3), // Templated
							// Inputs
							.reg_app_ecc_addr_protect_en(reg_app_ecc_addr_protect_en), // Templated
							.reg_app_ecc_bypass(reg_app_ecc_bypass), // Templated
							.reg_app_ecc_fault_detc_en(reg_app_ecc_fault_detc_en), // Templated
							.reg_app_pkt_crc_gen_dis(reg_app_pkt_crc_gen_dis), // Templated
							.reg_resv_pkt_match_lp_dt(reg_resv_pkt_match_lp_dt_pipe3[5:0]), // Templated
							.reg_resv_pkt_match_lp_dt_en(reg_resv_pkt_match_lp_dt_en_pipe3), // Templated
							.reg_sram_lcrc_err_oen(reg_sram_lcrc_err_oen[3]), // Templated
							.reg_video_fifo_empty_depend_cnt_mux(reg_video_fifo_empty_depend_cnt_mux), // Templated
							.clk_1M		(clk_1M),	 // Templated
							.fifo_wrclk	(fifo_wrclk3),	 // Templated
							.fifo_wrclk_rst_n(fifo_wrclk_rst_n3), // Templated
							.fifo_rdclk	(fifo_rdclk3),	 // Templated
							.fifo_rdclk_rst_n(fifo_rdclk_rst_n3), // Templated
							.in_csi_data	(pipe3_csi_data[(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0]), // Templated
							.in_bytes_en	(pipe3_bytes_en[(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0]), // Templated
							.in_header_en	(pipe3_header_en), // Templated
							.in_data_en	(pipe3_data_en), // Templated
							.in_data_type	(pipe3_data_type[5:0]), // Templated
							.in_virtual_channel(pipe3_virtual_channel[1:0]), // Templated
							.in_virtual_channel_x(pipe3_virtual_channel_x[(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0]), // Templated
							.in_word_count	(pipe3_word_count[15:0]), // Templated
							.in_aggr_id	(pipe3_aggr_id[3:0]), // Templated
							.in_pkt_crc	(pipe3_pkt_crc[31:0]), // Templated
							.in_pkt_crc_en	(pipe3_pkt_crc_en), // Templated
							.up_state	(up_state_video_pipe3), // Templated
							.line_delay_en	(line_delay_en3), // Templated
							.video_loss_en	(video_loss_en3), // Templated
							.time_window	(time_window3[16:0]), // Templated
							.reg_dft_tpram_config(reg_dft_tpram_config[8:0]), // Templated
							.reg_dft_sync_tpram_config(reg_dft_sync_tpram_config[9:0]), // Templated
							.app_aggregation_bypass(app_aggregation_bypass), // Templated
							.reg_video_pipe_en(reg_video_pipe_en[3]), // Templated
							.reg_last_byte_header_down_mux(reg_last_byte_header_down_mux), // Templated
							.reg_clear_resv_pkt_cnt_lp_pf(reg_clear_resv_pkt_cnt_lp_pf_pipe3), // Templated
							.reg_clear_resv_pkt_cnt_lp_ph(reg_clear_resv_pkt_cnt_lp_ph_pipe3), // Templated
							.reg_clear_resv_pkt_cnt_sp_le(reg_clear_resv_pkt_cnt_sp_le_pipe3), // Templated
							.reg_clear_resv_pkt_cnt_sp_ls(reg_clear_resv_pkt_cnt_sp_ls_pipe3), // Templated
							.reg_clear_resv_pkt_cnt_sp_fe(reg_clear_resv_pkt_cnt_sp_fe_pipe3), // Templated
							.reg_clear_resv_pkt_cnt_sp_fs(reg_clear_resv_pkt_cnt_sp_fs_pipe3), // Templated
							.reg_clear_app_full_cnt_async_fifo(reg_clear_app_full_cnt_async_fifo_pipe3), // Templated
							.reg_clear_app_full_cnt_sync_fifo(reg_clear_app_full_cnt_sync_fifo_pipe3), // Templated
							.reg_app_wr_idi_data_continue(reg_app_wr_idi_data_continue), // Templated
							.reg_dbg_pkt_num_nonzero_threshold(reg_dbg_pkt_num_nonzero_threshold[15:0]), // Templated
							.reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold(reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold[15:0])); // Templated

as6d_app_video_pipe_lane    u4_as6d_app_video_pipe_lane(/*AUTOINST*/
							// Outputs
							.ack_pre	(ack_pre4),	 // Templated
							.video_data_afifo_ecc_fault(video_data_afifo_ecc_fault4), // Templated
							.video_data_fwft_fifo_ecc_fault(video_data_fwft_fifo_ecc_fault4), // Templated
							.video_data_afifo_single_err(video_data_afifo_single_err4), // Templated
							.video_data_afifo_double_err(video_data_afifo_double_err4), // Templated
							.video_data_afifo_ovf_int(video_data_afifo_ovf_int4), // Templated
							.video_data_afifo_udf_int(video_data_afifo_udf_int4), // Templated
							.video_data_afifo_prog_full(video_data_afifo_prog_full4), // Templated
							.video_data_afifo_empty(video_data_afifo_empty4), // Templated
							.video_data_afifo_full(video_data_afifo_full4), // Templated
							.video_data_afifo_prog_empty(video_data_afifo_prog_empty4), // Templated
							.video_data_fwft_fifo_single_err(video_data_fwft_fifo_single_err4), // Templated
							.video_data_fwft_fifo_double_err(video_data_fwft_fifo_double_err4), // Templated
							.video_data_fwft_fifo_ovf_int(video_data_fwft_fifo_ovf_int4), // Templated
							.video_data_fwft_fifo_udf_int(video_data_fwft_fifo_udf_int4), // Templated
							.video_data_fwft_fifo_prog_full(video_data_fwft_fifo_prog_full4), // Templated
							.video_data_fwft_fifo_empty(video_data_fwft_fifo_empty4), // Templated
							.video_data_fwft_fifo_full(video_data_fwft_fifo_full4), // Templated
							.video_data_vld	(video_data_vld4), // Templated
							.video_data	(video_data4[(VIDEO_DATA_SIZE-1):0]), // Templated
							.ack		(ack4),		 // Templated
							.line_end	(line_end4),	 // Templated
							.video_loss	(video_loss4),	 // Templated
							.video_lock	(video_lock4),	 // Templated
							.fifo_rd_ctrl_cs(fifo_rd_ctrl_cs4[2:0]), // Templated
							.fs_detect_pipe	(fs_detect_pipe4), // Templated
							.fs_cnt_pipe	(fs_cnt_pipe4[15:0]), // Templated
							.empty_vld_aggregator0(empty_vld_pipe4_aggregator0), // Templated
							.empty_vld_aggregator1(empty_vld_pipe4_aggregator1), // Templated
							.empty_vld_aggregator2(empty_vld_pipe4_aggregator2), // Templated
							.empty_vld_aggregator3(empty_vld_pipe4_aggregator3), // Templated
							.ack_vld_aggregator0(ack_vld_pipe4_aggregator0), // Templated
							.ack_vld_aggregator1(ack_vld_pipe4_aggregator1), // Templated
							.ack_vld_aggregator2(ack_vld_pipe4_aggregator2), // Templated
							.ack_vld_aggregator3(ack_vld_pipe4_aggregator3), // Templated
							.line_end_vld_aggregator0(line_end_vld_pipe4_aggregator0), // Templated
							.line_end_vld_aggregator1(line_end_vld_pipe4_aggregator1), // Templated
							.line_end_vld_aggregator2(line_end_vld_pipe4_aggregator2), // Templated
							.line_end_vld_aggregator3(line_end_vld_pipe4_aggregator3), // Templated
							.video_pipe_data_aggre_bypass(video_pipe4_data_aggre_bypass[139:0]), // Templated
							.video_pipe_vld_aggre_bypass(video_pipe4_vld_aggre_bypass), // Templated
							.reg_rd_resv_pkt_cnt_lp_pf(reg_rd_resv_pkt_cnt_lp_pf_pipe4[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_lp_ph(reg_rd_resv_pkt_cnt_lp_ph_pipe4[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_le(reg_rd_resv_pkt_cnt_sp_le_pipe4[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_ls(reg_rd_resv_pkt_cnt_sp_ls_pipe4[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fe(reg_rd_resv_pkt_cnt_sp_fe_pipe4[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fs(reg_rd_resv_pkt_cnt_sp_fs_pipe4[31:0]), // Templated
							.reg_rd_app_full_cnt_sync_fifo(reg_rd_app_full_cnt_sync_fifo_pipe4[31:0]), // Templated
							.reg_rd_app_full_cnt_async_fifo(reg_rd_app_full_cnt_async_fifo_pipe4[31:0]), // Templated
							.reg_rd_dispatched_cnt_ready_for_sch(reg_rd_pipe4_dispatched_cnt_ready_for_sch[31:0]), // Templated
							.lcrc_err	(lcrc_err4),	 // Templated
							.reg_rd_dbg_pkt_num_nonzero_threshold_err(reg_rd_dbg_pkt_num_nonzero_threshold_err[4]), // Templated
							.reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err(reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err[4]), // Templated
							.video_pipe_date_type_for_concat_align(video_pipe_date_type_for_concat_align4[5:0]), // Templated
							.video_pipe_date_type_for_concat_align_vld(video_pipe_date_type_for_concat_align_vld4), // Templated
							// Inputs
							.reg_app_ecc_addr_protect_en(reg_app_ecc_addr_protect_en), // Templated
							.reg_app_ecc_bypass(reg_app_ecc_bypass), // Templated
							.reg_app_ecc_fault_detc_en(reg_app_ecc_fault_detc_en), // Templated
							.reg_app_pkt_crc_gen_dis(reg_app_pkt_crc_gen_dis), // Templated
							.reg_resv_pkt_match_lp_dt(reg_resv_pkt_match_lp_dt_pipe4[5:0]), // Templated
							.reg_resv_pkt_match_lp_dt_en(reg_resv_pkt_match_lp_dt_en_pipe4), // Templated
							.reg_sram_lcrc_err_oen(reg_sram_lcrc_err_oen[4]), // Templated
							.reg_video_fifo_empty_depend_cnt_mux(reg_video_fifo_empty_depend_cnt_mux), // Templated
							.clk_1M		(clk_1M),	 // Templated
							.fifo_wrclk	(fifo_wrclk4),	 // Templated
							.fifo_wrclk_rst_n(fifo_wrclk_rst_n4), // Templated
							.fifo_rdclk	(fifo_rdclk4),	 // Templated
							.fifo_rdclk_rst_n(fifo_rdclk_rst_n4), // Templated
							.in_csi_data	(pipe4_csi_data[(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0]), // Templated
							.in_bytes_en	(pipe4_bytes_en[(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0]), // Templated
							.in_header_en	(pipe4_header_en), // Templated
							.in_data_en	(pipe4_data_en), // Templated
							.in_data_type	(pipe4_data_type[5:0]), // Templated
							.in_virtual_channel(pipe4_virtual_channel[1:0]), // Templated
							.in_virtual_channel_x(pipe4_virtual_channel_x[(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0]), // Templated
							.in_word_count	(pipe4_word_count[15:0]), // Templated
							.in_aggr_id	(pipe4_aggr_id[3:0]), // Templated
							.in_pkt_crc	(pipe4_pkt_crc[31:0]), // Templated
							.in_pkt_crc_en	(pipe4_pkt_crc_en), // Templated
							.up_state	(up_state_video_pipe4), // Templated
							.line_delay_en	(line_delay_en4), // Templated
							.video_loss_en	(video_loss_en4), // Templated
							.time_window	(time_window4[16:0]), // Templated
							.reg_dft_tpram_config(reg_dft_tpram_config[8:0]), // Templated
							.reg_dft_sync_tpram_config(reg_dft_sync_tpram_config[9:0]), // Templated
							.app_aggregation_bypass(app_aggregation_bypass), // Templated
							.reg_video_pipe_en(reg_video_pipe_en[4]), // Templated
							.reg_last_byte_header_down_mux(reg_last_byte_header_down_mux), // Templated
							.reg_clear_resv_pkt_cnt_lp_pf(reg_clear_resv_pkt_cnt_lp_pf_pipe4), // Templated
							.reg_clear_resv_pkt_cnt_lp_ph(reg_clear_resv_pkt_cnt_lp_ph_pipe4), // Templated
							.reg_clear_resv_pkt_cnt_sp_le(reg_clear_resv_pkt_cnt_sp_le_pipe4), // Templated
							.reg_clear_resv_pkt_cnt_sp_ls(reg_clear_resv_pkt_cnt_sp_ls_pipe4), // Templated
							.reg_clear_resv_pkt_cnt_sp_fe(reg_clear_resv_pkt_cnt_sp_fe_pipe4), // Templated
							.reg_clear_resv_pkt_cnt_sp_fs(reg_clear_resv_pkt_cnt_sp_fs_pipe4), // Templated
							.reg_clear_app_full_cnt_async_fifo(reg_clear_app_full_cnt_async_fifo_pipe4), // Templated
							.reg_clear_app_full_cnt_sync_fifo(reg_clear_app_full_cnt_sync_fifo_pipe4), // Templated
							.reg_app_wr_idi_data_continue(reg_app_wr_idi_data_continue), // Templated
							.reg_dbg_pkt_num_nonzero_threshold(reg_dbg_pkt_num_nonzero_threshold[15:0]), // Templated
							.reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold(reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold[15:0])); // Templated
as6d_app_video_pipe_lane    u5_as6d_app_video_pipe_lane(/*AUTOINST*/
							// Outputs
							.ack_pre	(ack_pre5),	 // Templated
							.video_data_afifo_ecc_fault(video_data_afifo_ecc_fault5), // Templated
							.video_data_fwft_fifo_ecc_fault(video_data_fwft_fifo_ecc_fault5), // Templated
							.video_data_afifo_single_err(video_data_afifo_single_err5), // Templated
							.video_data_afifo_double_err(video_data_afifo_double_err5), // Templated
							.video_data_afifo_ovf_int(video_data_afifo_ovf_int5), // Templated
							.video_data_afifo_udf_int(video_data_afifo_udf_int5), // Templated
							.video_data_afifo_prog_full(video_data_afifo_prog_full5), // Templated
							.video_data_afifo_empty(video_data_afifo_empty5), // Templated
							.video_data_afifo_full(video_data_afifo_full5), // Templated
							.video_data_afifo_prog_empty(video_data_afifo_prog_empty5), // Templated
							.video_data_fwft_fifo_single_err(video_data_fwft_fifo_single_err5), // Templated
							.video_data_fwft_fifo_double_err(video_data_fwft_fifo_double_err5), // Templated
							.video_data_fwft_fifo_ovf_int(video_data_fwft_fifo_ovf_int5), // Templated
							.video_data_fwft_fifo_udf_int(video_data_fwft_fifo_udf_int5), // Templated
							.video_data_fwft_fifo_prog_full(video_data_fwft_fifo_prog_full5), // Templated
							.video_data_fwft_fifo_empty(video_data_fwft_fifo_empty5), // Templated
							.video_data_fwft_fifo_full(video_data_fwft_fifo_full5), // Templated
							.video_data_vld	(video_data_vld5), // Templated
							.video_data	(video_data5[(VIDEO_DATA_SIZE-1):0]), // Templated
							.ack		(ack5),		 // Templated
							.line_end	(line_end5),	 // Templated
							.video_loss	(video_loss5),	 // Templated
							.video_lock	(video_lock5),	 // Templated
							.fifo_rd_ctrl_cs(fifo_rd_ctrl_cs5[2:0]), // Templated
							.fs_detect_pipe	(fs_detect_pipe5), // Templated
							.fs_cnt_pipe	(fs_cnt_pipe5[15:0]), // Templated
							.empty_vld_aggregator0(empty_vld_pipe5_aggregator0), // Templated
							.empty_vld_aggregator1(empty_vld_pipe5_aggregator1), // Templated
							.empty_vld_aggregator2(empty_vld_pipe5_aggregator2), // Templated
							.empty_vld_aggregator3(empty_vld_pipe5_aggregator3), // Templated
							.ack_vld_aggregator0(ack_vld_pipe5_aggregator0), // Templated
							.ack_vld_aggregator1(ack_vld_pipe5_aggregator1), // Templated
							.ack_vld_aggregator2(ack_vld_pipe5_aggregator2), // Templated
							.ack_vld_aggregator3(ack_vld_pipe5_aggregator3), // Templated
							.line_end_vld_aggregator0(line_end_vld_pipe5_aggregator0), // Templated
							.line_end_vld_aggregator1(line_end_vld_pipe5_aggregator1), // Templated
							.line_end_vld_aggregator2(line_end_vld_pipe5_aggregator2), // Templated
							.line_end_vld_aggregator3(line_end_vld_pipe5_aggregator3), // Templated
							.video_pipe_data_aggre_bypass(video_pipe5_data_aggre_bypass[139:0]), // Templated
							.video_pipe_vld_aggre_bypass(video_pipe5_vld_aggre_bypass), // Templated
							.reg_rd_resv_pkt_cnt_lp_pf(reg_rd_resv_pkt_cnt_lp_pf_pipe5[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_lp_ph(reg_rd_resv_pkt_cnt_lp_ph_pipe5[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_le(reg_rd_resv_pkt_cnt_sp_le_pipe5[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_ls(reg_rd_resv_pkt_cnt_sp_ls_pipe5[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fe(reg_rd_resv_pkt_cnt_sp_fe_pipe5[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fs(reg_rd_resv_pkt_cnt_sp_fs_pipe5[31:0]), // Templated
							.reg_rd_app_full_cnt_sync_fifo(reg_rd_app_full_cnt_sync_fifo_pipe5[31:0]), // Templated
							.reg_rd_app_full_cnt_async_fifo(reg_rd_app_full_cnt_async_fifo_pipe5[31:0]), // Templated
							.reg_rd_dispatched_cnt_ready_for_sch(reg_rd_pipe5_dispatched_cnt_ready_for_sch[31:0]), // Templated
							.lcrc_err	(lcrc_err5),	 // Templated
							.reg_rd_dbg_pkt_num_nonzero_threshold_err(reg_rd_dbg_pkt_num_nonzero_threshold_err[5]), // Templated
							.reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err(reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err[5]), // Templated
							.video_pipe_date_type_for_concat_align(video_pipe_date_type_for_concat_align5[5:0]), // Templated
							.video_pipe_date_type_for_concat_align_vld(video_pipe_date_type_for_concat_align_vld5), // Templated
							// Inputs
							.reg_app_ecc_addr_protect_en(reg_app_ecc_addr_protect_en), // Templated
							.reg_app_ecc_bypass(reg_app_ecc_bypass), // Templated
							.reg_app_ecc_fault_detc_en(reg_app_ecc_fault_detc_en), // Templated
							.reg_app_pkt_crc_gen_dis(reg_app_pkt_crc_gen_dis), // Templated
							.reg_resv_pkt_match_lp_dt(reg_resv_pkt_match_lp_dt_pipe5[5:0]), // Templated
							.reg_resv_pkt_match_lp_dt_en(reg_resv_pkt_match_lp_dt_en_pipe5), // Templated
							.reg_sram_lcrc_err_oen(reg_sram_lcrc_err_oen[5]), // Templated
							.reg_video_fifo_empty_depend_cnt_mux(reg_video_fifo_empty_depend_cnt_mux), // Templated
							.clk_1M		(clk_1M),	 // Templated
							.fifo_wrclk	(fifo_wrclk5),	 // Templated
							.fifo_wrclk_rst_n(fifo_wrclk_rst_n5), // Templated
							.fifo_rdclk	(fifo_rdclk5),	 // Templated
							.fifo_rdclk_rst_n(fifo_rdclk_rst_n5), // Templated
							.in_csi_data	(pipe5_csi_data[(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0]), // Templated
							.in_bytes_en	(pipe5_bytes_en[(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0]), // Templated
							.in_header_en	(pipe5_header_en), // Templated
							.in_data_en	(pipe5_data_en), // Templated
							.in_data_type	(pipe5_data_type[5:0]), // Templated
							.in_virtual_channel(pipe5_virtual_channel[1:0]), // Templated
							.in_virtual_channel_x(pipe5_virtual_channel_x[(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0]), // Templated
							.in_word_count	(pipe5_word_count[15:0]), // Templated
							.in_aggr_id	(pipe5_aggr_id[3:0]), // Templated
							.in_pkt_crc	(pipe5_pkt_crc[31:0]), // Templated
							.in_pkt_crc_en	(pipe5_pkt_crc_en), // Templated
							.up_state	(up_state_video_pipe5), // Templated
							.line_delay_en	(line_delay_en5), // Templated
							.video_loss_en	(video_loss_en5), // Templated
							.time_window	(time_window5[16:0]), // Templated
							.reg_dft_tpram_config(reg_dft_tpram_config[8:0]), // Templated
							.reg_dft_sync_tpram_config(reg_dft_sync_tpram_config[9:0]), // Templated
							.app_aggregation_bypass(app_aggregation_bypass), // Templated
							.reg_video_pipe_en(reg_video_pipe_en[5]), // Templated
							.reg_last_byte_header_down_mux(reg_last_byte_header_down_mux), // Templated
							.reg_clear_resv_pkt_cnt_lp_pf(reg_clear_resv_pkt_cnt_lp_pf_pipe5), // Templated
							.reg_clear_resv_pkt_cnt_lp_ph(reg_clear_resv_pkt_cnt_lp_ph_pipe5), // Templated
							.reg_clear_resv_pkt_cnt_sp_le(reg_clear_resv_pkt_cnt_sp_le_pipe5), // Templated
							.reg_clear_resv_pkt_cnt_sp_ls(reg_clear_resv_pkt_cnt_sp_ls_pipe5), // Templated
							.reg_clear_resv_pkt_cnt_sp_fe(reg_clear_resv_pkt_cnt_sp_fe_pipe5), // Templated
							.reg_clear_resv_pkt_cnt_sp_fs(reg_clear_resv_pkt_cnt_sp_fs_pipe5), // Templated
							.reg_clear_app_full_cnt_async_fifo(reg_clear_app_full_cnt_async_fifo_pipe5), // Templated
							.reg_clear_app_full_cnt_sync_fifo(reg_clear_app_full_cnt_sync_fifo_pipe5), // Templated
							.reg_app_wr_idi_data_continue(reg_app_wr_idi_data_continue), // Templated
							.reg_dbg_pkt_num_nonzero_threshold(reg_dbg_pkt_num_nonzero_threshold[15:0]), // Templated
							.reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold(reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold[15:0])); // Templated
as6d_app_video_pipe_lane    u6_as6d_app_video_pipe_lane(/*AUTOINST*/
							// Outputs
							.ack_pre	(ack_pre6),	 // Templated
							.video_data_afifo_ecc_fault(video_data_afifo_ecc_fault6), // Templated
							.video_data_fwft_fifo_ecc_fault(video_data_fwft_fifo_ecc_fault6), // Templated
							.video_data_afifo_single_err(video_data_afifo_single_err6), // Templated
							.video_data_afifo_double_err(video_data_afifo_double_err6), // Templated
							.video_data_afifo_ovf_int(video_data_afifo_ovf_int6), // Templated
							.video_data_afifo_udf_int(video_data_afifo_udf_int6), // Templated
							.video_data_afifo_prog_full(video_data_afifo_prog_full6), // Templated
							.video_data_afifo_empty(video_data_afifo_empty6), // Templated
							.video_data_afifo_full(video_data_afifo_full6), // Templated
							.video_data_afifo_prog_empty(video_data_afifo_prog_empty6), // Templated
							.video_data_fwft_fifo_single_err(video_data_fwft_fifo_single_err6), // Templated
							.video_data_fwft_fifo_double_err(video_data_fwft_fifo_double_err6), // Templated
							.video_data_fwft_fifo_ovf_int(video_data_fwft_fifo_ovf_int6), // Templated
							.video_data_fwft_fifo_udf_int(video_data_fwft_fifo_udf_int6), // Templated
							.video_data_fwft_fifo_prog_full(video_data_fwft_fifo_prog_full6), // Templated
							.video_data_fwft_fifo_empty(video_data_fwft_fifo_empty6), // Templated
							.video_data_fwft_fifo_full(video_data_fwft_fifo_full6), // Templated
							.video_data_vld	(video_data_vld6), // Templated
							.video_data	(video_data6[(VIDEO_DATA_SIZE-1):0]), // Templated
							.ack		(ack6),		 // Templated
							.line_end	(line_end6),	 // Templated
							.video_loss	(video_loss6),	 // Templated
							.video_lock	(video_lock6),	 // Templated
							.fifo_rd_ctrl_cs(fifo_rd_ctrl_cs6[2:0]), // Templated
							.fs_detect_pipe	(fs_detect_pipe6), // Templated
							.fs_cnt_pipe	(fs_cnt_pipe6[15:0]), // Templated
							.empty_vld_aggregator0(empty_vld_pipe6_aggregator0), // Templated
							.empty_vld_aggregator1(empty_vld_pipe6_aggregator1), // Templated
							.empty_vld_aggregator2(empty_vld_pipe6_aggregator2), // Templated
							.empty_vld_aggregator3(empty_vld_pipe6_aggregator3), // Templated
							.ack_vld_aggregator0(ack_vld_pipe6_aggregator0), // Templated
							.ack_vld_aggregator1(ack_vld_pipe6_aggregator1), // Templated
							.ack_vld_aggregator2(ack_vld_pipe6_aggregator2), // Templated
							.ack_vld_aggregator3(ack_vld_pipe6_aggregator3), // Templated
							.line_end_vld_aggregator0(line_end_vld_pipe6_aggregator0), // Templated
							.line_end_vld_aggregator1(line_end_vld_pipe6_aggregator1), // Templated
							.line_end_vld_aggregator2(line_end_vld_pipe6_aggregator2), // Templated
							.line_end_vld_aggregator3(line_end_vld_pipe6_aggregator3), // Templated
							.video_pipe_data_aggre_bypass(video_pipe6_data_aggre_bypass[139:0]), // Templated
							.video_pipe_vld_aggre_bypass(video_pipe6_vld_aggre_bypass), // Templated
							.reg_rd_resv_pkt_cnt_lp_pf(reg_rd_resv_pkt_cnt_lp_pf_pipe6[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_lp_ph(reg_rd_resv_pkt_cnt_lp_ph_pipe6[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_le(reg_rd_resv_pkt_cnt_sp_le_pipe6[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_ls(reg_rd_resv_pkt_cnt_sp_ls_pipe6[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fe(reg_rd_resv_pkt_cnt_sp_fe_pipe6[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fs(reg_rd_resv_pkt_cnt_sp_fs_pipe6[31:0]), // Templated
							.reg_rd_app_full_cnt_sync_fifo(reg_rd_app_full_cnt_sync_fifo_pipe6[31:0]), // Templated
							.reg_rd_app_full_cnt_async_fifo(reg_rd_app_full_cnt_async_fifo_pipe6[31:0]), // Templated
							.reg_rd_dispatched_cnt_ready_for_sch(reg_rd_pipe6_dispatched_cnt_ready_for_sch[31:0]), // Templated
							.lcrc_err	(lcrc_err6),	 // Templated
							.reg_rd_dbg_pkt_num_nonzero_threshold_err(reg_rd_dbg_pkt_num_nonzero_threshold_err[6]), // Templated
							.reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err(reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err[6]), // Templated
							.video_pipe_date_type_for_concat_align(video_pipe_date_type_for_concat_align6[5:0]), // Templated
							.video_pipe_date_type_for_concat_align_vld(video_pipe_date_type_for_concat_align_vld6), // Templated
							// Inputs
							.reg_app_ecc_addr_protect_en(reg_app_ecc_addr_protect_en), // Templated
							.reg_app_ecc_bypass(reg_app_ecc_bypass), // Templated
							.reg_app_ecc_fault_detc_en(reg_app_ecc_fault_detc_en), // Templated
							.reg_app_pkt_crc_gen_dis(reg_app_pkt_crc_gen_dis), // Templated
							.reg_resv_pkt_match_lp_dt(reg_resv_pkt_match_lp_dt_pipe6[5:0]), // Templated
							.reg_resv_pkt_match_lp_dt_en(reg_resv_pkt_match_lp_dt_en_pipe6), // Templated
							.reg_sram_lcrc_err_oen(reg_sram_lcrc_err_oen[6]), // Templated
							.reg_video_fifo_empty_depend_cnt_mux(reg_video_fifo_empty_depend_cnt_mux), // Templated
							.clk_1M		(clk_1M),	 // Templated
							.fifo_wrclk	(fifo_wrclk6),	 // Templated
							.fifo_wrclk_rst_n(fifo_wrclk_rst_n6), // Templated
							.fifo_rdclk	(fifo_rdclk6),	 // Templated
							.fifo_rdclk_rst_n(fifo_rdclk_rst_n6), // Templated
							.in_csi_data	(pipe6_csi_data[(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0]), // Templated
							.in_bytes_en	(pipe6_bytes_en[(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0]), // Templated
							.in_header_en	(pipe6_header_en), // Templated
							.in_data_en	(pipe6_data_en), // Templated
							.in_data_type	(pipe6_data_type[5:0]), // Templated
							.in_virtual_channel(pipe6_virtual_channel[1:0]), // Templated
							.in_virtual_channel_x(pipe6_virtual_channel_x[(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0]), // Templated
							.in_word_count	(pipe6_word_count[15:0]), // Templated
							.in_aggr_id	(pipe6_aggr_id[3:0]), // Templated
							.in_pkt_crc	(pipe6_pkt_crc[31:0]), // Templated
							.in_pkt_crc_en	(pipe6_pkt_crc_en), // Templated
							.up_state	(up_state_video_pipe6), // Templated
							.line_delay_en	(line_delay_en6), // Templated
							.video_loss_en	(video_loss_en6), // Templated
							.time_window	(time_window6[16:0]), // Templated
							.reg_dft_tpram_config(reg_dft_tpram_config[8:0]), // Templated
							.reg_dft_sync_tpram_config(reg_dft_sync_tpram_config[9:0]), // Templated
							.app_aggregation_bypass(app_aggregation_bypass), // Templated
							.reg_video_pipe_en(reg_video_pipe_en[6]), // Templated
							.reg_last_byte_header_down_mux(reg_last_byte_header_down_mux), // Templated
							.reg_clear_resv_pkt_cnt_lp_pf(reg_clear_resv_pkt_cnt_lp_pf_pipe6), // Templated
							.reg_clear_resv_pkt_cnt_lp_ph(reg_clear_resv_pkt_cnt_lp_ph_pipe6), // Templated
							.reg_clear_resv_pkt_cnt_sp_le(reg_clear_resv_pkt_cnt_sp_le_pipe6), // Templated
							.reg_clear_resv_pkt_cnt_sp_ls(reg_clear_resv_pkt_cnt_sp_ls_pipe6), // Templated
							.reg_clear_resv_pkt_cnt_sp_fe(reg_clear_resv_pkt_cnt_sp_fe_pipe6), // Templated
							.reg_clear_resv_pkt_cnt_sp_fs(reg_clear_resv_pkt_cnt_sp_fs_pipe6), // Templated
							.reg_clear_app_full_cnt_async_fifo(reg_clear_app_full_cnt_async_fifo_pipe6), // Templated
							.reg_clear_app_full_cnt_sync_fifo(reg_clear_app_full_cnt_sync_fifo_pipe6), // Templated
							.reg_app_wr_idi_data_continue(reg_app_wr_idi_data_continue), // Templated
							.reg_dbg_pkt_num_nonzero_threshold(reg_dbg_pkt_num_nonzero_threshold[15:0]), // Templated
							.reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold(reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold[15:0])); // Templated
as6d_app_video_pipe_lane    u7_as6d_app_video_pipe_lane(/*AUTOINST*/
							// Outputs
							.ack_pre	(ack_pre7),	 // Templated
							.video_data_afifo_ecc_fault(video_data_afifo_ecc_fault7), // Templated
							.video_data_fwft_fifo_ecc_fault(video_data_fwft_fifo_ecc_fault7), // Templated
							.video_data_afifo_single_err(video_data_afifo_single_err7), // Templated
							.video_data_afifo_double_err(video_data_afifo_double_err7), // Templated
							.video_data_afifo_ovf_int(video_data_afifo_ovf_int7), // Templated
							.video_data_afifo_udf_int(video_data_afifo_udf_int7), // Templated
							.video_data_afifo_prog_full(video_data_afifo_prog_full7), // Templated
							.video_data_afifo_empty(video_data_afifo_empty7), // Templated
							.video_data_afifo_full(video_data_afifo_full7), // Templated
							.video_data_afifo_prog_empty(video_data_afifo_prog_empty7), // Templated
							.video_data_fwft_fifo_single_err(video_data_fwft_fifo_single_err7), // Templated
							.video_data_fwft_fifo_double_err(video_data_fwft_fifo_double_err7), // Templated
							.video_data_fwft_fifo_ovf_int(video_data_fwft_fifo_ovf_int7), // Templated
							.video_data_fwft_fifo_udf_int(video_data_fwft_fifo_udf_int7), // Templated
							.video_data_fwft_fifo_prog_full(video_data_fwft_fifo_prog_full7), // Templated
							.video_data_fwft_fifo_empty(video_data_fwft_fifo_empty7), // Templated
							.video_data_fwft_fifo_full(video_data_fwft_fifo_full7), // Templated
							.video_data_vld	(video_data_vld7), // Templated
							.video_data	(video_data7[(VIDEO_DATA_SIZE-1):0]), // Templated
							.ack		(ack7),		 // Templated
							.line_end	(line_end7),	 // Templated
							.video_loss	(video_loss7),	 // Templated
							.video_lock	(video_lock7),	 // Templated
							.fifo_rd_ctrl_cs(fifo_rd_ctrl_cs7[2:0]), // Templated
							.fs_detect_pipe	(fs_detect_pipe7), // Templated
							.fs_cnt_pipe	(fs_cnt_pipe7[15:0]), // Templated
							.empty_vld_aggregator0(empty_vld_pipe7_aggregator0), // Templated
							.empty_vld_aggregator1(empty_vld_pipe7_aggregator1), // Templated
							.empty_vld_aggregator2(empty_vld_pipe7_aggregator2), // Templated
							.empty_vld_aggregator3(empty_vld_pipe7_aggregator3), // Templated
							.ack_vld_aggregator0(ack_vld_pipe7_aggregator0), // Templated
							.ack_vld_aggregator1(ack_vld_pipe7_aggregator1), // Templated
							.ack_vld_aggregator2(ack_vld_pipe7_aggregator2), // Templated
							.ack_vld_aggregator3(ack_vld_pipe7_aggregator3), // Templated
							.line_end_vld_aggregator0(line_end_vld_pipe7_aggregator0), // Templated
							.line_end_vld_aggregator1(line_end_vld_pipe7_aggregator1), // Templated
							.line_end_vld_aggregator2(line_end_vld_pipe7_aggregator2), // Templated
							.line_end_vld_aggregator3(line_end_vld_pipe7_aggregator3), // Templated
							.video_pipe_data_aggre_bypass(video_pipe7_data_aggre_bypass[139:0]), // Templated
							.video_pipe_vld_aggre_bypass(video_pipe7_vld_aggre_bypass), // Templated
							.reg_rd_resv_pkt_cnt_lp_pf(reg_rd_resv_pkt_cnt_lp_pf_pipe7[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_lp_ph(reg_rd_resv_pkt_cnt_lp_ph_pipe7[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_le(reg_rd_resv_pkt_cnt_sp_le_pipe7[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_ls(reg_rd_resv_pkt_cnt_sp_ls_pipe7[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fe(reg_rd_resv_pkt_cnt_sp_fe_pipe7[31:0]), // Templated
							.reg_rd_resv_pkt_cnt_sp_fs(reg_rd_resv_pkt_cnt_sp_fs_pipe7[31:0]), // Templated
							.reg_rd_app_full_cnt_sync_fifo(reg_rd_app_full_cnt_sync_fifo_pipe7[31:0]), // Templated
							.reg_rd_app_full_cnt_async_fifo(reg_rd_app_full_cnt_async_fifo_pipe7[31:0]), // Templated
							.reg_rd_dispatched_cnt_ready_for_sch(reg_rd_pipe7_dispatched_cnt_ready_for_sch[31:0]), // Templated
							.lcrc_err	(lcrc_err7),	 // Templated
							.reg_rd_dbg_pkt_num_nonzero_threshold_err(reg_rd_dbg_pkt_num_nonzero_threshold_err[7]), // Templated
							.reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err(reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err[7]), // Templated
							.video_pipe_date_type_for_concat_align(video_pipe_date_type_for_concat_align7[5:0]), // Templated
							.video_pipe_date_type_for_concat_align_vld(video_pipe_date_type_for_concat_align_vld7), // Templated
							// Inputs
							.reg_app_ecc_addr_protect_en(reg_app_ecc_addr_protect_en), // Templated
							.reg_app_ecc_bypass(reg_app_ecc_bypass), // Templated
							.reg_app_ecc_fault_detc_en(reg_app_ecc_fault_detc_en), // Templated
							.reg_app_pkt_crc_gen_dis(reg_app_pkt_crc_gen_dis), // Templated
							.reg_resv_pkt_match_lp_dt(reg_resv_pkt_match_lp_dt_pipe7[5:0]), // Templated
							.reg_resv_pkt_match_lp_dt_en(reg_resv_pkt_match_lp_dt_en_pipe7), // Templated
							.reg_sram_lcrc_err_oen(reg_sram_lcrc_err_oen[7]), // Templated
							.reg_video_fifo_empty_depend_cnt_mux(reg_video_fifo_empty_depend_cnt_mux), // Templated
							.clk_1M		(clk_1M),	 // Templated
							.fifo_wrclk	(fifo_wrclk7),	 // Templated
							.fifo_wrclk_rst_n(fifo_wrclk_rst_n7), // Templated
							.fifo_rdclk	(fifo_rdclk7),	 // Templated
							.fifo_rdclk_rst_n(fifo_rdclk_rst_n7), // Templated
							.in_csi_data	(pipe7_csi_data[(`MEP_CSI2_DEVICE_IDI_CSIDATA_SIZE-1):0]), // Templated
							.in_bytes_en	(pipe7_bytes_en[(`MEP_CSI2_DEVICE_IDI_DATA_BYTEEN_WIDTH-1):0]), // Templated
							.in_header_en	(pipe7_header_en), // Templated
							.in_data_en	(pipe7_data_en), // Templated
							.in_data_type	(pipe7_data_type[5:0]), // Templated
							.in_virtual_channel(pipe7_virtual_channel[1:0]), // Templated
							.in_virtual_channel_x(pipe7_virtual_channel_x[(`MEP_CSI2_DEVICE_VCX_DWIDTH-1):0]), // Templated
							.in_word_count	(pipe7_word_count[15:0]), // Templated
							.in_aggr_id	(pipe7_aggr_id[3:0]), // Templated
							.in_pkt_crc	(pipe7_pkt_crc[31:0]), // Templated
							.in_pkt_crc_en	(pipe7_pkt_crc_en), // Templated
							.up_state	(up_state_video_pipe7), // Templated
							.line_delay_en	(line_delay_en7), // Templated
							.video_loss_en	(video_loss_en7), // Templated
							.time_window	(time_window7[16:0]), // Templated
							.reg_dft_tpram_config(reg_dft_tpram_config[8:0]), // Templated
							.reg_dft_sync_tpram_config(reg_dft_sync_tpram_config[9:0]), // Templated
							.app_aggregation_bypass(app_aggregation_bypass), // Templated
							.reg_video_pipe_en(reg_video_pipe_en[7]), // Templated
							.reg_last_byte_header_down_mux(reg_last_byte_header_down_mux), // Templated
							.reg_clear_resv_pkt_cnt_lp_pf(reg_clear_resv_pkt_cnt_lp_pf_pipe7), // Templated
							.reg_clear_resv_pkt_cnt_lp_ph(reg_clear_resv_pkt_cnt_lp_ph_pipe7), // Templated
							.reg_clear_resv_pkt_cnt_sp_le(reg_clear_resv_pkt_cnt_sp_le_pipe7), // Templated
							.reg_clear_resv_pkt_cnt_sp_ls(reg_clear_resv_pkt_cnt_sp_ls_pipe7), // Templated
							.reg_clear_resv_pkt_cnt_sp_fe(reg_clear_resv_pkt_cnt_sp_fe_pipe7), // Templated
							.reg_clear_resv_pkt_cnt_sp_fs(reg_clear_resv_pkt_cnt_sp_fs_pipe7), // Templated
							.reg_clear_app_full_cnt_async_fifo(reg_clear_app_full_cnt_async_fifo_pipe7), // Templated
							.reg_clear_app_full_cnt_sync_fifo(reg_clear_app_full_cnt_sync_fifo_pipe7), // Templated
							.reg_app_wr_idi_data_continue(reg_app_wr_idi_data_continue), // Templated
							.reg_dbg_pkt_num_nonzero_threshold(reg_dbg_pkt_num_nonzero_threshold[15:0]), // Templated
							.reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold(reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold[15:0])); // Templated

                            
assign fifo_rdclk          =   {fifo_rdclk7,
                                fifo_rdclk6,  
                                fifo_rdclk5,
                                fifo_rdclk4,
                                fifo_rdclk3,
                                fifo_rdclk2,  
                                fifo_rdclk1,
                                fifo_rdclk0};
                            
assign fifo_rdclk_rst_n    =   {fifo_rdclk_rst_n7,
                                fifo_rdclk_rst_n6,  
                                fifo_rdclk_rst_n5,
                                fifo_rdclk_rst_n4,
                                fifo_rdclk_rst_n3,
                                fifo_rdclk_rst_n2,  
                                fifo_rdclk_rst_n1,
                                fifo_rdclk_rst_n0};

assign pipe_fifo_full_pre  =   {video_data_fwft_fifo_full7,
                                video_data_fwft_fifo_full6,
                                video_data_fwft_fifo_full5,
                                video_data_fwft_fifo_full4,
                                video_data_fwft_fifo_full3,
                                video_data_fwft_fifo_full2,
                                video_data_fwft_fifo_full1,
                                video_data_fwft_fifo_full0};

generate for(j=0;j<=7;j=j+1)begin:pulse_cnt_pipe_fifo_bk
    as6d_app_pulse_cnt#(
        .CNT_WDTH(1)
    ) as6d_app_pulse_cnt_pipe_fifo(
        .cnt    (reg_rd_pipe_fifo_full[j]),    
        .clk    (fifo_rdclk[j]),    
        .rst_n  (fifo_rdclk_rst_n[j]),    
        .clear  (pipe_fifo_full_clear[j]),  
        .pulse  (pipe_fifo_full_pre[j])    
    );
end
endgenerate


endmodule
