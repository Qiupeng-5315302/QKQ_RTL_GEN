
package idi_vip_pkg

    `include "/data/proj/as6t28d/wa/xuhaiqiang/my_tb/idi_bus_vip/idi_interface.sv"
    `include "/data/proj/as6t28d/wa/xuhaiqiang/my_tb/idi_bus_vip/idi_config.sv"
    `include "/data/proj/as6t28d/wa/xuhaiqiang/my_tb/idi_bus_vip/idi_driver.sv"
    `include "/data/proj/as6t28d/wa/xuhaiqiang/my_tb/idi_bus_vip/idi_monitor.sv"
    `include "/data/proj/as6t28d/wa/xuhaiqiang/my_tb/idi_bus_vip/idi_env.sv"

endpackage : idi_vip_pkg
