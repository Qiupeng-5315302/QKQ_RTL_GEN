
`include "as6d_app_all_includes.vh"
module as6d_app_lcrc_check(/*AUTOARG*/
   // Outputs
   out_data_vld, out_data, out_crc_err,
   // Inputs
   clk, rst_n, in_data_vld, in_data, in_crc_vld, in_crc
   );
    //inputs
    input               								clk;
    input               								rst_n;
    input                                               in_data_vld;
    input      [139:0]                                  in_data;
    input              								    in_crc_vld;
    input      [31:0]									in_crc;

    //outputs
    output                                              out_data_vld;
    output     [139:0]                                  out_data;
    output                                              out_crc_err;

    //signal definition
    localparam              PACKET_HEADER = 4'b0001;
    localparam              PACKET_DATA   = 2'b10;
    localparam              PACKET_FOOTER = 2'b10;
    wire        [31:0]      crc_32_out;
    reg         [31:0]      crc_32_reg;
    wire                    sob_in;
    wire                    eob_in;
    reg         [139:0]     data_in_d1;
    reg         [139:0]     data_in_d2;
    reg         [31:0]      crc_in_d1;
    reg         [31:0]      crc_in_d2;
    reg                     data_vld_in_d1;
    reg                     data_vld_in_d2;
    reg                     crc_vld_in_d1;
    reg                     crc_vld_in_d2;
    reg                     sob_in_d1;
    reg                     eob_in_d1;
    reg         [31:0]      di;
    reg         [31:0]      crc;
    reg         [139:0]     out_data;
    reg                     out_data_vld;
    reg                     out_crc_err;
    reg         [3:0]       data_in_d1_lock_high_4bit;

    //logic body
    assign sob_in  =   in_data_vld & (in_data[135:132] == PACKET_HEADER);
    assign eob_in  =   in_data_vld & (in_data[133:132] == PACKET_FOOTER);

    always@(posedge clk or negedge rst_n)begin
        if(!rst_n)begin
            data_in_d1 <= 140'd0;
            data_in_d2 <= 140'd0;
            crc_in_d1  <= 32'd0;
            crc_in_d2  <= 32'd0;
        end
        else begin
            data_in_d1 <= in_data;
            data_in_d2 <= data_in_d1;
            crc_in_d1  <= in_crc;
            crc_in_d2  <= crc_in_d1;
        end
    end

    always@(posedge clk or negedge rst_n)begin
        if(!rst_n)begin
            data_vld_in_d1 <= 1'd0;
            data_vld_in_d2 <= 1'd0;
            crc_vld_in_d1  <= 1'd0;
            crc_vld_in_d2  <= 1'd0;
            sob_in_d1      <= 1'd0;
            eob_in_d1      <= 1'd0;
        end
        else begin
            data_vld_in_d1 <= in_data_vld;
            data_vld_in_d2 <= data_vld_in_d1;
            crc_vld_in_d1  <= in_crc_vld;
            crc_vld_in_d2  <= crc_vld_in_d1;
            sob_in_d1      <= sob_in;
            eob_in_d1      <= eob_in;
        end
    end

    always @(posedge clk or negedge rst_n)begin
        if(!rst_n)begin
            di <= 32'b0;
        end
        else if(in_data_vld)begin
            di <= next_din_140(in_data);
        end
    end
    
    always@(posedge clk or negedge rst_n)begin
        if(!rst_n)
            crc <= 32'd0;
        else if(data_vld_in_d1)begin
            if(sob_in_d1)begin
                crc <= next_crc_140(di,32'd0);
            end
            else begin
                crc <= next_crc_140(di,crc);
            end
        end
    end

    always@(posedge clk or negedge rst_n)begin
        if(!rst_n)
            data_in_d1_lock_high_4bit <= 4'd0;
        else if(data_vld_in_d1)begin
            if(eob_in_d1)begin
                data_in_d1_lock_high_4bit <= data_in_d1[139:136];
            end
        end
    end

    always@(posedge clk or negedge rst_n)begin
        if(!rst_n)begin
            out_data     <= 140'd0;
            out_data_vld <= 1'd0;
        end
        else if(data_vld_in_d2)begin
            out_data     <= data_in_d2;
            out_data_vld <= 1'd1;
        end
        else if(crc_vld_in_d2)begin
            out_data     <= {data_in_d1_lock_high_4bit,4'd0,crc,100'd0};
            out_data_vld <= 1'd1;
        end
        else begin
            out_data_vld <= 1'd0;
        end
    end

    always@(posedge clk or negedge rst_n)begin
        if(!rst_n)begin
            out_crc_err <= 1'b0;
        end
        else if(crc_vld_in_d2)begin
            out_crc_err <= |(crc_in_d2 ^ crc);
        end
        else begin
            out_crc_err <= 1'b0;
        end
    end

    function automatic [31:0] next_din_140;
        input [139:0]  d;
        reg [31:0]  next_d;
        begin
            next_d[31] = d[ 5] ^d[ 8] ^d[ 9] ^d[11] ^d[15] ^d[23] ^d[24] ^d[25] ^d[27] ^d[28] ^d[29] ^d[30] ^d[31] ^d[33] ^d[36] ^d[43] ^d[44] ^d[46] ^d[47] ^d[49] ^d[52] ^d[53] ^d[54] ^d[57] ^d[59] ^d[60] ^d[62] ^d[64] ^d[65] ^d[66] ^d[67] ^d[71] ^d[72] ^d[78] ^d[80] ^d[81] ^d[82] ^d[83] ^d[84] ^d[86] ^d[93] ^d[94] ^d[95] ^d[96] ^d[97] ^d[98] ^d[100] ^d[102] ^d[103] ^d[105] ^d[109] ^d[110] ^d[112] ^d[113] ^d[115] ^d[116] ^d[117] ^d[118] ^d[122] ^d[124] ^d[125] ^d[126] ^d[127] ^d[131] ^d[133] ^d[134] ^d[135] ^d[136] ;
            next_d[30] = d[ 4] ^d[ 7] ^d[ 8] ^d[10] ^d[14] ^d[22] ^d[23] ^d[24] ^d[26] ^d[27] ^d[28] ^d[29] ^d[30] ^d[32] ^d[35] ^d[42] ^d[43] ^d[45] ^d[46] ^d[48] ^d[51] ^d[52] ^d[53] ^d[56] ^d[58] ^d[59] ^d[61] ^d[63] ^d[64] ^d[65] ^d[66] ^d[70] ^d[71] ^d[77] ^d[79] ^d[80] ^d[81] ^d[82] ^d[83] ^d[85] ^d[92] ^d[93] ^d[94] ^d[95] ^d[96] ^d[97] ^d[99] ^d[101] ^d[102] ^d[104] ^d[108] ^d[109] ^d[111] ^d[112] ^d[114] ^d[115] ^d[116] ^d[117] ^d[121] ^d[123] ^d[124] ^d[125] ^d[126] ^d[130] ^d[132] ^d[133] ^d[134] ^d[135] ;
            next_d[29] = d[ 3] ^d[ 6] ^d[ 7] ^d[ 9] ^d[13] ^d[21] ^d[22] ^d[23] ^d[25] ^d[26] ^d[27] ^d[28] ^d[29] ^d[31] ^d[34] ^d[41] ^d[42] ^d[44] ^d[45] ^d[47] ^d[50] ^d[51] ^d[52] ^d[55] ^d[57] ^d[58] ^d[60] ^d[62] ^d[63] ^d[64] ^d[65] ^d[69] ^d[70] ^d[76] ^d[78] ^d[79] ^d[80] ^d[81] ^d[82] ^d[84] ^d[91] ^d[92] ^d[93] ^d[94] ^d[95] ^d[96] ^d[98] ^d[100] ^d[101] ^d[103] ^d[107] ^d[108] ^d[110] ^d[111] ^d[113] ^d[114] ^d[115] ^d[116] ^d[120] ^d[122] ^d[123] ^d[124] ^d[125] ^d[129] ^d[131] ^d[132] ^d[133] ^d[134] ;
            next_d[28] = d[ 2] ^d[ 5] ^d[ 6] ^d[ 8] ^d[12] ^d[20] ^d[21] ^d[22] ^d[24] ^d[25] ^d[26] ^d[27] ^d[28] ^d[30] ^d[33] ^d[40] ^d[41] ^d[43] ^d[44] ^d[46] ^d[49] ^d[50] ^d[51] ^d[54] ^d[56] ^d[57] ^d[59] ^d[61] ^d[62] ^d[63] ^d[64] ^d[68] ^d[69] ^d[75] ^d[77] ^d[78] ^d[79] ^d[80] ^d[81] ^d[83] ^d[90] ^d[91] ^d[92] ^d[93] ^d[94] ^d[95] ^d[97] ^d[99] ^d[100] ^d[102] ^d[106] ^d[107] ^d[109] ^d[110] ^d[112] ^d[113] ^d[114] ^d[115] ^d[119] ^d[121] ^d[122] ^d[123] ^d[124] ^d[128] ^d[130] ^d[131] ^d[132] ^d[133] ^d[139] ;
            next_d[27] = d[ 1] ^d[ 4] ^d[ 5] ^d[ 7] ^d[11] ^d[19] ^d[20] ^d[21] ^d[23] ^d[24] ^d[25] ^d[26] ^d[27] ^d[29] ^d[32] ^d[39] ^d[40] ^d[42] ^d[43] ^d[45] ^d[48] ^d[49] ^d[50] ^d[53] ^d[55] ^d[56] ^d[58] ^d[60] ^d[61] ^d[62] ^d[63] ^d[67] ^d[68] ^d[74] ^d[76] ^d[77] ^d[78] ^d[79] ^d[80] ^d[82] ^d[89] ^d[90] ^d[91] ^d[92] ^d[93] ^d[94] ^d[96] ^d[98] ^d[99] ^d[101] ^d[105] ^d[106] ^d[108] ^d[109] ^d[111] ^d[112] ^d[113] ^d[114] ^d[118] ^d[120] ^d[121] ^d[122] ^d[123] ^d[127] ^d[129] ^d[130] ^d[131] ^d[132] ^d[138] ^d[139] ;
            next_d[26] = d[ 0] ^d[ 3] ^d[ 4] ^d[ 6] ^d[10] ^d[18] ^d[19] ^d[20] ^d[22] ^d[23] ^d[24] ^d[25] ^d[26] ^d[28] ^d[31] ^d[38] ^d[39] ^d[41] ^d[42] ^d[44] ^d[47] ^d[48] ^d[49] ^d[52] ^d[54] ^d[55] ^d[57] ^d[59] ^d[60] ^d[61] ^d[62] ^d[66] ^d[67] ^d[73] ^d[75] ^d[76] ^d[77] ^d[78] ^d[79] ^d[81] ^d[88] ^d[89] ^d[90] ^d[91] ^d[92] ^d[93] ^d[95] ^d[97] ^d[98] ^d[100] ^d[104] ^d[105] ^d[107] ^d[108] ^d[110] ^d[111] ^d[112] ^d[113] ^d[117] ^d[119] ^d[120] ^d[121] ^d[122] ^d[126] ^d[128] ^d[129] ^d[130] ^d[131] ^d[137] ^d[138] ;
            next_d[25] = d[ 2] ^d[ 3] ^d[ 8] ^d[11] ^d[15] ^d[17] ^d[18] ^d[19] ^d[21] ^d[22] ^d[28] ^d[29] ^d[31] ^d[33] ^d[36] ^d[37] ^d[38] ^d[40] ^d[41] ^d[44] ^d[48] ^d[49] ^d[51] ^d[52] ^d[56] ^d[57] ^d[58] ^d[61] ^d[62] ^d[64] ^d[67] ^d[71] ^d[74] ^d[75] ^d[76] ^d[77] ^d[81] ^d[82] ^d[83] ^d[84] ^d[86] ^d[87] ^d[88] ^d[89] ^d[90] ^d[91] ^d[92] ^d[93] ^d[95] ^d[98] ^d[99] ^d[100] ^d[102] ^d[104] ^d[105] ^d[106] ^d[107] ^d[111] ^d[113] ^d[115] ^d[117] ^d[119] ^d[120] ^d[121] ^d[122] ^d[124] ^d[126] ^d[128] ^d[129] ^d[130] ^d[131] ^d[133] ^d[134] ^d[135] ^d[137] ;
            next_d[24] = d[ 1] ^d[ 2] ^d[ 7] ^d[10] ^d[14] ^d[16] ^d[17] ^d[18] ^d[20] ^d[21] ^d[27] ^d[28] ^d[30] ^d[32] ^d[35] ^d[36] ^d[37] ^d[39] ^d[40] ^d[43] ^d[47] ^d[48] ^d[50] ^d[51] ^d[55] ^d[56] ^d[57] ^d[60] ^d[61] ^d[63] ^d[66] ^d[70] ^d[73] ^d[74] ^d[75] ^d[76] ^d[80] ^d[81] ^d[82] ^d[83] ^d[85] ^d[86] ^d[87] ^d[88] ^d[89] ^d[90] ^d[91] ^d[92] ^d[94] ^d[97] ^d[98] ^d[99] ^d[101] ^d[103] ^d[104] ^d[105] ^d[106] ^d[110] ^d[112] ^d[114] ^d[116] ^d[118] ^d[119] ^d[120] ^d[121] ^d[123] ^d[125] ^d[127] ^d[128] ^d[129] ^d[130] ^d[132] ^d[133] ^d[134] ^d[136] ;
            next_d[23] = d[ 0] ^d[ 1] ^d[ 6] ^d[ 9] ^d[13] ^d[15] ^d[16] ^d[17] ^d[19] ^d[20] ^d[26] ^d[27] ^d[29] ^d[31] ^d[34] ^d[35] ^d[36] ^d[38] ^d[39] ^d[42] ^d[46] ^d[47] ^d[49] ^d[50] ^d[54] ^d[55] ^d[56] ^d[59] ^d[60] ^d[62] ^d[65] ^d[69] ^d[72] ^d[73] ^d[74] ^d[75] ^d[79] ^d[80] ^d[81] ^d[82] ^d[84] ^d[85] ^d[86] ^d[87] ^d[88] ^d[89] ^d[90] ^d[91] ^d[93] ^d[96] ^d[97] ^d[98] ^d[100] ^d[102] ^d[103] ^d[104] ^d[105] ^d[109] ^d[111] ^d[113] ^d[115] ^d[117] ^d[118] ^d[119] ^d[120] ^d[122] ^d[124] ^d[126] ^d[127] ^d[128] ^d[129] ^d[131] ^d[132] ^d[133] ^d[135] ;
            next_d[22] = d[ 0] ^d[ 9] ^d[11] ^d[12] ^d[14] ^d[16] ^d[18] ^d[19] ^d[23] ^d[24] ^d[26] ^d[27] ^d[29] ^d[31] ^d[34] ^d[35] ^d[36] ^d[37] ^d[38] ^d[41] ^d[43] ^d[44] ^d[45] ^d[47] ^d[48] ^d[52] ^d[55] ^d[57] ^d[58] ^d[60] ^d[61] ^d[62] ^d[65] ^d[66] ^d[67] ^d[68] ^d[73] ^d[74] ^d[79] ^d[82] ^d[85] ^d[87] ^d[88] ^d[89] ^d[90] ^d[92] ^d[93] ^d[94] ^d[98] ^d[99] ^d[100] ^d[101] ^d[104] ^d[105] ^d[108] ^d[109] ^d[113] ^d[114] ^d[115] ^d[119] ^d[121] ^d[122] ^d[123] ^d[124] ^d[128] ^d[130] ^d[132] ^d[133] ^d[135] ^d[136] ;
            next_d[21] = d[ 5] ^d[ 9] ^d[10] ^d[13] ^d[17] ^d[18] ^d[22] ^d[24] ^d[26] ^d[27] ^d[29] ^d[31] ^d[34] ^d[35] ^d[37] ^d[40] ^d[42] ^d[49] ^d[51] ^d[52] ^d[53] ^d[56] ^d[61] ^d[62] ^d[71] ^d[73] ^d[80] ^d[82] ^d[83] ^d[87] ^d[88] ^d[89] ^d[91] ^d[92] ^d[94] ^d[95] ^d[96] ^d[99] ^d[102] ^d[104] ^d[105] ^d[107] ^d[108] ^d[109] ^d[110] ^d[114] ^d[115] ^d[116] ^d[117] ^d[120] ^d[121] ^d[123] ^d[124] ^d[125] ^d[126] ^d[129] ^d[132] ^d[133] ^d[136] ^d[139] ;
            next_d[20] = d[ 4] ^d[ 8] ^d[ 9] ^d[12] ^d[16] ^d[17] ^d[21] ^d[23] ^d[25] ^d[26] ^d[28] ^d[30] ^d[33] ^d[34] ^d[36] ^d[39] ^d[41] ^d[48] ^d[50] ^d[51] ^d[52] ^d[55] ^d[60] ^d[61] ^d[70] ^d[72] ^d[79] ^d[81] ^d[82] ^d[86] ^d[87] ^d[88] ^d[90] ^d[91] ^d[93] ^d[94] ^d[95] ^d[98] ^d[101] ^d[103] ^d[104] ^d[106] ^d[107] ^d[108] ^d[109] ^d[113] ^d[114] ^d[115] ^d[116] ^d[119] ^d[120] ^d[122] ^d[123] ^d[124] ^d[125] ^d[128] ^d[131] ^d[132] ^d[135] ^d[138] ^d[139] ;
            next_d[19] = d[ 3] ^d[ 7] ^d[ 8] ^d[11] ^d[15] ^d[16] ^d[20] ^d[22] ^d[24] ^d[25] ^d[27] ^d[29] ^d[32] ^d[33] ^d[35] ^d[38] ^d[40] ^d[47] ^d[49] ^d[50] ^d[51] ^d[54] ^d[59] ^d[60] ^d[69] ^d[71] ^d[78] ^d[80] ^d[81] ^d[85] ^d[86] ^d[87] ^d[89] ^d[90] ^d[92] ^d[93] ^d[94] ^d[97] ^d[100] ^d[102] ^d[103] ^d[105] ^d[106] ^d[107] ^d[108] ^d[112] ^d[113] ^d[114] ^d[115] ^d[118] ^d[119] ^d[121] ^d[122] ^d[123] ^d[124] ^d[127] ^d[130] ^d[131] ^d[134] ^d[137] ^d[138] ^d[139] ;
            next_d[18] = d[ 2] ^d[ 6] ^d[ 7] ^d[10] ^d[14] ^d[15] ^d[19] ^d[21] ^d[23] ^d[24] ^d[26] ^d[28] ^d[31] ^d[32] ^d[34] ^d[37] ^d[39] ^d[46] ^d[48] ^d[49] ^d[50] ^d[53] ^d[58] ^d[59] ^d[68] ^d[70] ^d[77] ^d[79] ^d[80] ^d[84] ^d[85] ^d[86] ^d[88] ^d[89] ^d[91] ^d[92] ^d[93] ^d[96] ^d[99] ^d[101] ^d[102] ^d[104] ^d[105] ^d[106] ^d[107] ^d[111] ^d[112] ^d[113] ^d[114] ^d[117] ^d[118] ^d[120] ^d[121] ^d[122] ^d[123] ^d[126] ^d[129] ^d[130] ^d[133] ^d[136] ^d[137] ^d[138] ;
            next_d[17] = d[ 1] ^d[ 5] ^d[ 6] ^d[ 9] ^d[13] ^d[14] ^d[18] ^d[20] ^d[22] ^d[23] ^d[25] ^d[27] ^d[30] ^d[31] ^d[33] ^d[36] ^d[38] ^d[45] ^d[47] ^d[48] ^d[49] ^d[52] ^d[57] ^d[58] ^d[67] ^d[69] ^d[76] ^d[78] ^d[79] ^d[83] ^d[84] ^d[85] ^d[87] ^d[88] ^d[90] ^d[91] ^d[92] ^d[95] ^d[98] ^d[100] ^d[101] ^d[103] ^d[104] ^d[105] ^d[106] ^d[110] ^d[111] ^d[112] ^d[113] ^d[116] ^d[117] ^d[119] ^d[120] ^d[121] ^d[122] ^d[125] ^d[128] ^d[129] ^d[132] ^d[135] ^d[136] ^d[137] ^d[139] ;
            next_d[16] = d[ 0] ^d[ 4] ^d[ 5] ^d[ 8] ^d[12] ^d[13] ^d[17] ^d[19] ^d[21] ^d[22] ^d[24] ^d[26] ^d[29] ^d[30] ^d[32] ^d[35] ^d[37] ^d[44] ^d[46] ^d[47] ^d[48] ^d[51] ^d[56] ^d[57] ^d[66] ^d[68] ^d[75] ^d[77] ^d[78] ^d[82] ^d[83] ^d[84] ^d[86] ^d[87] ^d[89] ^d[90] ^d[91] ^d[94] ^d[97] ^d[99] ^d[100] ^d[102] ^d[103] ^d[104] ^d[105] ^d[109] ^d[110] ^d[111] ^d[112] ^d[115] ^d[116] ^d[118] ^d[119] ^d[120] ^d[121] ^d[124] ^d[127] ^d[128] ^d[131] ^d[134] ^d[135] ^d[136] ^d[138] ;
            next_d[15] = d[ 3] ^d[ 4] ^d[ 5] ^d[ 7] ^d[ 8] ^d[ 9] ^d[12] ^d[15] ^d[16] ^d[18] ^d[20] ^d[21] ^d[24] ^d[27] ^d[30] ^d[33] ^d[34] ^d[44] ^d[45] ^d[49] ^d[50] ^d[52] ^d[53] ^d[54] ^d[55] ^d[56] ^d[57] ^d[59] ^d[60] ^d[62] ^d[64] ^d[66] ^d[71] ^d[72] ^d[74] ^d[76] ^d[77] ^d[78] ^d[80] ^d[84] ^d[85] ^d[88] ^d[89] ^d[90] ^d[94] ^d[95] ^d[97] ^d[99] ^d[100] ^d[101] ^d[104] ^d[105] ^d[108] ^d[111] ^d[112] ^d[113] ^d[114] ^d[116] ^d[119] ^d[120] ^d[122] ^d[123] ^d[124] ^d[125] ^d[130] ^d[131] ^d[136] ^d[137] ^d[139] ;
            next_d[14] = d[ 2] ^d[ 3] ^d[ 4] ^d[ 6] ^d[ 7] ^d[ 8] ^d[11] ^d[14] ^d[15] ^d[17] ^d[19] ^d[20] ^d[23] ^d[26] ^d[29] ^d[32] ^d[33] ^d[43] ^d[44] ^d[48] ^d[49] ^d[51] ^d[52] ^d[53] ^d[54] ^d[55] ^d[56] ^d[58] ^d[59] ^d[61] ^d[63] ^d[65] ^d[70] ^d[71] ^d[73] ^d[75] ^d[76] ^d[77] ^d[79] ^d[83] ^d[84] ^d[87] ^d[88] ^d[89] ^d[93] ^d[94] ^d[96] ^d[98] ^d[99] ^d[100] ^d[103] ^d[104] ^d[107] ^d[110] ^d[111] ^d[112] ^d[113] ^d[115] ^d[118] ^d[119] ^d[121] ^d[122] ^d[123] ^d[124] ^d[129] ^d[130] ^d[135] ^d[136] ^d[138] ^d[139] ;
            next_d[13] = d[ 1] ^d[ 2] ^d[ 3] ^d[ 5] ^d[ 6] ^d[ 7] ^d[10] ^d[13] ^d[14] ^d[16] ^d[18] ^d[19] ^d[22] ^d[25] ^d[28] ^d[31] ^d[32] ^d[42] ^d[43] ^d[47] ^d[48] ^d[50] ^d[51] ^d[52] ^d[53] ^d[54] ^d[55] ^d[57] ^d[58] ^d[60] ^d[62] ^d[64] ^d[69] ^d[70] ^d[72] ^d[74] ^d[75] ^d[76] ^d[78] ^d[82] ^d[83] ^d[86] ^d[87] ^d[88] ^d[92] ^d[93] ^d[95] ^d[97] ^d[98] ^d[99] ^d[102] ^d[103] ^d[106] ^d[109] ^d[110] ^d[111] ^d[112] ^d[114] ^d[117] ^d[118] ^d[120] ^d[121] ^d[122] ^d[123] ^d[128] ^d[129] ^d[134] ^d[135] ^d[137] ^d[138] ;
            next_d[12] = d[ 0] ^d[ 1] ^d[ 2] ^d[ 4] ^d[ 5] ^d[ 6] ^d[ 9] ^d[12] ^d[13] ^d[15] ^d[17] ^d[18] ^d[21] ^d[24] ^d[27] ^d[30] ^d[31] ^d[41] ^d[42] ^d[46] ^d[47] ^d[49] ^d[50] ^d[51] ^d[52] ^d[53] ^d[54] ^d[56] ^d[57] ^d[59] ^d[61] ^d[63] ^d[68] ^d[69] ^d[71] ^d[73] ^d[74] ^d[75] ^d[77] ^d[81] ^d[82] ^d[85] ^d[86] ^d[87] ^d[91] ^d[92] ^d[94] ^d[96] ^d[97] ^d[98] ^d[101] ^d[102] ^d[105] ^d[108] ^d[109] ^d[110] ^d[111] ^d[113] ^d[116] ^d[117] ^d[119] ^d[120] ^d[121] ^d[122] ^d[127] ^d[128] ^d[133] ^d[134] ^d[136] ^d[137] ;
            next_d[11] = d[ 0] ^d[ 1] ^d[ 3] ^d[ 4] ^d[ 9] ^d[12] ^d[14] ^d[15] ^d[16] ^d[17] ^d[20] ^d[24] ^d[25] ^d[26] ^d[27] ^d[28] ^d[31] ^d[33] ^d[36] ^d[40] ^d[41] ^d[43] ^d[44] ^d[45] ^d[47] ^d[48] ^d[50] ^d[51] ^d[54] ^d[55] ^d[56] ^d[57] ^d[58] ^d[59] ^d[64] ^d[65] ^d[66] ^d[68] ^d[70] ^d[71] ^d[73] ^d[74] ^d[76] ^d[78] ^d[82] ^d[83] ^d[85] ^d[90] ^d[91] ^d[94] ^d[98] ^d[101] ^d[102] ^d[103] ^d[104] ^d[105] ^d[107] ^d[108] ^d[113] ^d[117] ^d[119] ^d[120] ^d[121] ^d[122] ^d[124] ^d[125] ^d[131] ^d[132] ^d[134] ;
            next_d[10] = d[ 0] ^d[ 2] ^d[ 3] ^d[ 5] ^d[ 9] ^d[13] ^d[14] ^d[16] ^d[19] ^d[26] ^d[28] ^d[29] ^d[31] ^d[32] ^d[33] ^d[35] ^d[36] ^d[39] ^d[40] ^d[42] ^d[50] ^d[52] ^d[55] ^d[56] ^d[58] ^d[59] ^d[60] ^d[62] ^d[63] ^d[66] ^d[69] ^d[70] ^d[71] ^d[73] ^d[75] ^d[77] ^d[78] ^d[80] ^d[83] ^d[86] ^d[89] ^d[90] ^d[94] ^d[95] ^d[96] ^d[98] ^d[101] ^d[104] ^d[105] ^d[106] ^d[107] ^d[109] ^d[110] ^d[113] ^d[115] ^d[117] ^d[119] ^d[120] ^d[121] ^d[122] ^d[123] ^d[125] ^d[126] ^d[127] ^d[130] ^d[134] ^d[135] ^d[136] ^d[139] ;
            next_d[ 9] = d[ 1] ^d[ 2] ^d[ 4] ^d[ 5] ^d[ 9] ^d[11] ^d[12] ^d[13] ^d[18] ^d[23] ^d[24] ^d[29] ^d[32] ^d[33] ^d[34] ^d[35] ^d[36] ^d[38] ^d[39] ^d[41] ^d[43] ^d[44] ^d[46] ^d[47] ^d[51] ^d[52] ^d[53] ^d[55] ^d[58] ^d[60] ^d[61] ^d[64] ^d[66] ^d[67] ^d[68] ^d[69] ^d[70] ^d[71] ^d[74] ^d[76] ^d[77] ^d[78] ^d[79] ^d[80] ^d[81] ^d[83] ^d[84] ^d[85] ^d[86] ^d[88] ^d[89] ^d[96] ^d[98] ^d[102] ^d[104] ^d[106] ^d[108] ^d[110] ^d[113] ^d[114] ^d[115] ^d[117] ^d[119] ^d[120] ^d[121] ^d[127] ^d[129] ^d[131] ^d[136] ^d[138] ;
            next_d[ 8] = d[ 0] ^d[ 1] ^d[ 3] ^d[ 4] ^d[ 8] ^d[10] ^d[11] ^d[12] ^d[17] ^d[22] ^d[23] ^d[28] ^d[31] ^d[32] ^d[33] ^d[34] ^d[35] ^d[37] ^d[38] ^d[40] ^d[42] ^d[43] ^d[45] ^d[46] ^d[50] ^d[51] ^d[52] ^d[54] ^d[57] ^d[59] ^d[60] ^d[63] ^d[65] ^d[66] ^d[67] ^d[68] ^d[69] ^d[70] ^d[73] ^d[75] ^d[76] ^d[77] ^d[78] ^d[79] ^d[80] ^d[82] ^d[83] ^d[84] ^d[85] ^d[87] ^d[88] ^d[95] ^d[97] ^d[101] ^d[103] ^d[105] ^d[107] ^d[109] ^d[112] ^d[113] ^d[114] ^d[116] ^d[118] ^d[119] ^d[120] ^d[126] ^d[128] ^d[130] ^d[135] ^d[137] ^d[139] ;
            next_d[ 7] = d[ 0] ^d[ 2] ^d[ 3] ^d[ 5] ^d[ 7] ^d[ 8] ^d[10] ^d[15] ^d[16] ^d[21] ^d[22] ^d[23] ^d[24] ^d[25] ^d[28] ^d[29] ^d[32] ^d[34] ^d[37] ^d[39] ^d[41] ^d[42] ^d[43] ^d[45] ^d[46] ^d[47] ^d[50] ^d[51] ^d[52] ^d[54] ^d[56] ^d[57] ^d[58] ^d[60] ^d[68] ^d[69] ^d[71] ^d[74] ^d[75] ^d[76] ^d[77] ^d[79] ^d[80] ^d[87] ^d[93] ^d[95] ^d[97] ^d[98] ^d[103] ^d[104] ^d[105] ^d[106] ^d[108] ^d[109] ^d[110] ^d[111] ^d[116] ^d[119] ^d[122] ^d[124] ^d[126] ^d[129] ^d[131] ^d[133] ^d[135] ^d[138] ;
            next_d[ 6] = d[ 1] ^d[ 2] ^d[ 4] ^d[ 5] ^d[ 6] ^d[ 7] ^d[ 8] ^d[11] ^d[14] ^d[20] ^d[21] ^d[22] ^d[25] ^d[29] ^d[30] ^d[38] ^d[40] ^d[41] ^d[42] ^d[43] ^d[45] ^d[47] ^d[50] ^d[51] ^d[52] ^d[54] ^d[55] ^d[56] ^d[60] ^d[62] ^d[64] ^d[65] ^d[66] ^d[68] ^d[70] ^d[71] ^d[72] ^d[73] ^d[74] ^d[75] ^d[76] ^d[79] ^d[80] ^d[81] ^d[82] ^d[83] ^d[84] ^d[92] ^d[93] ^d[95] ^d[98] ^d[100] ^d[104] ^d[107] ^d[108] ^d[112] ^d[113] ^d[116] ^d[117] ^d[121] ^d[122] ^d[123] ^d[124] ^d[126] ^d[127] ^d[128] ^d[130] ^d[131] ^d[132] ^d[133] ^d[135] ^d[136] ^d[137] ^d[139] ;
            next_d[ 5] = d[ 0] ^d[ 1] ^d[ 3] ^d[ 4] ^d[ 5] ^d[ 6] ^d[ 7] ^d[10] ^d[13] ^d[19] ^d[20] ^d[21] ^d[24] ^d[28] ^d[29] ^d[37] ^d[39] ^d[40] ^d[41] ^d[42] ^d[44] ^d[46] ^d[49] ^d[50] ^d[51] ^d[53] ^d[54] ^d[55] ^d[59] ^d[61] ^d[63] ^d[64] ^d[65] ^d[67] ^d[69] ^d[70] ^d[71] ^d[72] ^d[73] ^d[74] ^d[75] ^d[78] ^d[79] ^d[80] ^d[81] ^d[82] ^d[83] ^d[91] ^d[92] ^d[94] ^d[97] ^d[99] ^d[103] ^d[106] ^d[107] ^d[111] ^d[112] ^d[115] ^d[116] ^d[120] ^d[121] ^d[122] ^d[123] ^d[125] ^d[126] ^d[127] ^d[129] ^d[130] ^d[131] ^d[132] ^d[134] ^d[135] ^d[136] ^d[138] ^d[139] ;
            next_d[ 4] = d[ 0] ^d[ 2] ^d[ 3] ^d[ 4] ^d[ 6] ^d[ 8] ^d[11] ^d[12] ^d[15] ^d[18] ^d[19] ^d[20] ^d[24] ^d[25] ^d[29] ^d[30] ^d[31] ^d[33] ^d[38] ^d[39] ^d[40] ^d[41] ^d[44] ^d[45] ^d[46] ^d[47] ^d[48] ^d[50] ^d[57] ^d[58] ^d[59] ^d[63] ^d[65] ^d[67] ^d[68] ^d[69] ^d[70] ^d[73] ^d[74] ^d[77] ^d[79] ^d[83] ^d[84] ^d[86] ^d[90] ^d[91] ^d[94] ^d[95] ^d[97] ^d[100] ^d[103] ^d[106] ^d[109] ^d[111] ^d[112] ^d[113] ^d[114] ^d[116] ^d[117] ^d[118] ^d[119] ^d[120] ^d[121] ^d[127] ^d[128] ^d[129] ^d[130] ^d[136] ^d[137] ^d[138] ^d[139] ;
            next_d[ 3] = d[ 1] ^d[ 2] ^d[ 3] ^d[ 7] ^d[ 8] ^d[ 9] ^d[10] ^d[14] ^d[15] ^d[17] ^d[18] ^d[19] ^d[25] ^d[27] ^d[31] ^d[32] ^d[33] ^d[36] ^d[37] ^d[38] ^d[39] ^d[40] ^d[45] ^d[52] ^d[53] ^d[54] ^d[56] ^d[58] ^d[59] ^d[60] ^d[65] ^d[68] ^d[69] ^d[71] ^d[73] ^d[76] ^d[80] ^d[81] ^d[84] ^d[85] ^d[86] ^d[89] ^d[90] ^d[95] ^d[97] ^d[98] ^d[99] ^d[100] ^d[103] ^d[108] ^d[109] ^d[111] ^d[119] ^d[120] ^d[122] ^d[124] ^d[125] ^d[128] ^d[129] ^d[131] ^d[133] ^d[134] ^d[137] ^d[138] ;
            next_d[ 2] = d[ 0] ^d[ 1] ^d[ 2] ^d[ 6] ^d[ 7] ^d[ 8] ^d[ 9] ^d[13] ^d[14] ^d[16] ^d[17] ^d[18] ^d[24] ^d[26] ^d[30] ^d[31] ^d[32] ^d[35] ^d[36] ^d[37] ^d[38] ^d[39] ^d[44] ^d[51] ^d[52] ^d[53] ^d[55] ^d[57] ^d[58] ^d[59] ^d[64] ^d[67] ^d[68] ^d[70] ^d[72] ^d[75] ^d[79] ^d[80] ^d[83] ^d[84] ^d[85] ^d[88] ^d[89] ^d[94] ^d[96] ^d[97] ^d[98] ^d[99] ^d[102] ^d[107] ^d[108] ^d[110] ^d[118] ^d[119] ^d[121] ^d[123] ^d[124] ^d[127] ^d[128] ^d[130] ^d[132] ^d[133] ^d[136] ^d[137] ^d[139] ;
            next_d[ 1] = d[ 0] ^d[ 1] ^d[ 6] ^d[ 7] ^d[ 9] ^d[11] ^d[12] ^d[13] ^d[16] ^d[17] ^d[24] ^d[27] ^d[28] ^d[33] ^d[34] ^d[35] ^d[37] ^d[38] ^d[44] ^d[46] ^d[47] ^d[49] ^d[50] ^d[51] ^d[53] ^d[56] ^d[58] ^d[59] ^d[60] ^d[62] ^d[63] ^d[64] ^d[65] ^d[69] ^d[72] ^d[74] ^d[79] ^d[80] ^d[81] ^d[86] ^d[87] ^d[88] ^d[94] ^d[100] ^d[101] ^d[102] ^d[103] ^d[105] ^d[106] ^d[107] ^d[110] ^d[112] ^d[113] ^d[115] ^d[116] ^d[120] ^d[123] ^d[124] ^d[125] ^d[129] ^d[132] ^d[133] ^d[134] ^d[138] ;
            next_d[ 0] = d[ 0] ^d[ 6] ^d[ 9] ^d[10] ^d[12] ^d[16] ^d[24] ^d[25] ^d[26] ^d[28] ^d[29] ^d[30] ^d[31] ^d[32] ^d[34] ^d[37] ^d[44] ^d[45] ^d[47] ^d[48] ^d[50] ^d[53] ^d[54] ^d[55] ^d[58] ^d[60] ^d[61] ^d[63] ^d[65] ^d[66] ^d[67] ^d[68] ^d[72] ^d[73] ^d[79] ^d[81] ^d[82] ^d[83] ^d[84] ^d[85] ^d[87] ^d[94] ^d[95] ^d[96] ^d[97] ^d[98] ^d[99] ^d[101] ^d[103] ^d[104] ^d[106] ^d[110] ^d[111] ^d[113] ^d[114] ^d[116] ^d[117] ^d[118] ^d[119] ^d[123] ^d[125] ^d[126] ^d[127] ^d[128] ^d[132] ^d[134] ^d[135] ^d[136] ^d[137] ;
            next_din_140 = next_d;
        end
    endfunction

    function automatic [31:0] next_crc_140;
        input [31:0]  d;
        input [31:0]  c;
        reg [31:0]  next_c;
        begin
            next_c[31] = d[31] ^c[28] ^c[27] ^c[26] ^c[25] ^c[23] ^c[19] ^c[18] ^c[17] ^c[16] ^c[14] ^c[10] ^c[ 9] ^c[ 8] ^c[ 7] ^c[ 5] ^c[ 4] ^c[ 2] ^c[ 1] ;
            next_c[30] = d[30] ^c[27] ^c[26] ^c[25] ^c[24] ^c[22] ^c[18] ^c[17] ^c[16] ^c[15] ^c[13] ^c[ 9] ^c[ 8] ^c[ 7] ^c[ 6] ^c[ 4] ^c[ 3] ^c[ 1] ^c[ 0] ;
            next_c[29] = d[29] ^c[26] ^c[25] ^c[24] ^c[23] ^c[21] ^c[17] ^c[16] ^c[15] ^c[14] ^c[12] ^c[ 8] ^c[ 7] ^c[ 6] ^c[ 5] ^c[ 3] ^c[ 2] ^c[ 0] ;
            next_c[28] = d[28] ^c[31] ^c[25] ^c[24] ^c[23] ^c[22] ^c[20] ^c[16] ^c[15] ^c[14] ^c[13] ^c[11] ^c[ 7] ^c[ 6] ^c[ 5] ^c[ 4] ^c[ 2] ^c[ 1] ;
            next_c[27] = d[27] ^c[31] ^c[30] ^c[24] ^c[23] ^c[22] ^c[21] ^c[19] ^c[15] ^c[14] ^c[13] ^c[12] ^c[10] ^c[ 6] ^c[ 5] ^c[ 4] ^c[ 3] ^c[ 1] ^c[ 0] ;
            next_c[26] = d[26] ^c[30] ^c[29] ^c[23] ^c[22] ^c[21] ^c[20] ^c[18] ^c[14] ^c[13] ^c[12] ^c[11] ^c[ 9] ^c[ 5] ^c[ 4] ^c[ 3] ^c[ 2] ^c[ 0] ;
            next_c[25] = d[25] ^c[29] ^c[27] ^c[26] ^c[25] ^c[23] ^c[22] ^c[21] ^c[20] ^c[18] ^c[16] ^c[14] ^c[13] ^c[12] ^c[11] ^c[ 9] ^c[ 7] ^c[ 5] ^c[ 3] ;
            next_c[24] = d[24] ^c[28] ^c[26] ^c[25] ^c[24] ^c[22] ^c[21] ^c[20] ^c[19] ^c[17] ^c[15] ^c[13] ^c[12] ^c[11] ^c[10] ^c[ 8] ^c[ 6] ^c[ 4] ^c[ 2] ;
            next_c[23] = d[23] ^c[27] ^c[25] ^c[24] ^c[23] ^c[21] ^c[20] ^c[19] ^c[18] ^c[16] ^c[14] ^c[12] ^c[11] ^c[10] ^c[ 9] ^c[ 7] ^c[ 5] ^c[ 3] ^c[ 1] ;
            next_c[22] = d[22] ^c[28] ^c[27] ^c[25] ^c[24] ^c[22] ^c[20] ^c[16] ^c[15] ^c[14] ^c[13] ^c[11] ^c[ 7] ^c[ 6] ^c[ 5] ^c[ 1] ^c[ 0] ;
            next_c[21] = d[21] ^c[31] ^c[28] ^c[25] ^c[24] ^c[21] ^c[18] ^c[17] ^c[16] ^c[15] ^c[13] ^c[12] ^c[ 9] ^c[ 8] ^c[ 7] ^c[ 6] ^c[ 2] ^c[ 1] ^c[ 0] ;
            next_c[20] = d[20] ^c[31] ^c[30] ^c[27] ^c[24] ^c[23] ^c[20] ^c[17] ^c[16] ^c[15] ^c[14] ^c[12] ^c[11] ^c[ 8] ^c[ 7] ^c[ 6] ^c[ 5] ^c[ 1] ^c[ 0] ;
            next_c[19] = d[19] ^c[31] ^c[30] ^c[29] ^c[26] ^c[23] ^c[22] ^c[19] ^c[16] ^c[15] ^c[14] ^c[13] ^c[11] ^c[10] ^c[ 7] ^c[ 6] ^c[ 5] ^c[ 4] ^c[ 0] ;
            next_c[18] = d[18] ^c[30] ^c[29] ^c[28] ^c[25] ^c[22] ^c[21] ^c[18] ^c[15] ^c[14] ^c[13] ^c[12] ^c[10] ^c[ 9] ^c[ 6] ^c[ 5] ^c[ 4] ^c[ 3] ;
            next_c[17] = d[17] ^c[31] ^c[29] ^c[28] ^c[27] ^c[24] ^c[21] ^c[20] ^c[17] ^c[14] ^c[13] ^c[12] ^c[11] ^c[ 9] ^c[ 8] ^c[ 5] ^c[ 4] ^c[ 3] ^c[ 2] ;
            next_c[16] = d[16] ^c[30] ^c[28] ^c[27] ^c[26] ^c[23] ^c[20] ^c[19] ^c[16] ^c[13] ^c[12] ^c[11] ^c[10] ^c[ 8] ^c[ 7] ^c[ 4] ^c[ 3] ^c[ 2] ^c[ 1] ;
            next_c[15] = d[15] ^c[31] ^c[29] ^c[28] ^c[23] ^c[22] ^c[17] ^c[16] ^c[15] ^c[14] ^c[12] ^c[11] ^c[ 8] ^c[ 6] ^c[ 5] ^c[ 4] ^c[ 3] ^c[ 0] ;
            next_c[14] = d[14] ^c[31] ^c[30] ^c[28] ^c[27] ^c[22] ^c[21] ^c[16] ^c[15] ^c[14] ^c[13] ^c[11] ^c[10] ^c[ 7] ^c[ 5] ^c[ 4] ^c[ 3] ^c[ 2] ;
            next_c[13] = d[13] ^c[30] ^c[29] ^c[27] ^c[26] ^c[21] ^c[20] ^c[15] ^c[14] ^c[13] ^c[12] ^c[10] ^c[ 9] ^c[ 6] ^c[ 4] ^c[ 3] ^c[ 2] ^c[ 1] ;
            next_c[12] = d[12] ^c[29] ^c[28] ^c[26] ^c[25] ^c[20] ^c[19] ^c[14] ^c[13] ^c[12] ^c[11] ^c[ 9] ^c[ 8] ^c[ 5] ^c[ 3] ^c[ 2] ^c[ 1] ^c[ 0] ;
            next_c[11] = d[11] ^c[26] ^c[24] ^c[23] ^c[17] ^c[16] ^c[14] ^c[13] ^c[12] ^c[11] ^c[ 9] ^c[ 5] ^c[ 0] ;
            next_c[10] = d[10] ^c[31] ^c[28] ^c[27] ^c[26] ^c[22] ^c[19] ^c[18] ^c[17] ^c[15] ^c[14] ^c[13] ^c[12] ^c[11] ^c[ 9] ^c[ 7] ^c[ 5] ^c[ 2] ^c[ 1] ;
            next_c[ 9] = d[ 9] ^c[30] ^c[28] ^c[23] ^c[21] ^c[19] ^c[13] ^c[12] ^c[11] ^c[ 9] ^c[ 7] ^c[ 6] ^c[ 5] ^c[ 2] ^c[ 0] ;
            next_c[ 8] = d[ 8] ^c[31] ^c[29] ^c[27] ^c[22] ^c[20] ^c[18] ^c[12] ^c[11] ^c[10] ^c[ 8] ^c[ 6] ^c[ 5] ^c[ 4] ^c[ 1] ;
            next_c[ 7] = d[ 7] ^c[30] ^c[27] ^c[25] ^c[23] ^c[21] ^c[18] ^c[16] ^c[14] ^c[11] ^c[ 8] ^c[ 3] ^c[ 2] ^c[ 1] ^c[ 0] ;
            next_c[ 6] = d[ 6] ^c[31] ^c[29] ^c[28] ^c[27] ^c[25] ^c[24] ^c[23] ^c[22] ^c[20] ^c[19] ^c[18] ^c[16] ^c[15] ^c[14] ^c[13] ^c[ 9] ^c[ 8] ^c[ 5] ^c[ 4] ^c[ 0] ;
            next_c[ 5] = d[ 5] ^c[31] ^c[30] ^c[28] ^c[27] ^c[26] ^c[24] ^c[23] ^c[22] ^c[21] ^c[19] ^c[18] ^c[17] ^c[15] ^c[14] ^c[13] ^c[12] ^c[ 8] ^c[ 7] ^c[ 4] ^c[ 3] ;
            next_c[ 4] = d[ 4] ^c[31] ^c[30] ^c[29] ^c[28] ^c[22] ^c[21] ^c[20] ^c[19] ^c[13] ^c[12] ^c[11] ^c[10] ^c[ 9] ^c[ 8] ^c[ 6] ^c[ 5] ^c[ 4] ^c[ 3] ^c[ 1] ;
            next_c[ 3] = d[ 3] ^c[30] ^c[29] ^c[26] ^c[25] ^c[23] ^c[21] ^c[20] ^c[17] ^c[16] ^c[14] ^c[12] ^c[11] ^c[ 3] ^c[ 1] ^c[ 0] ;
            next_c[ 2] = d[ 2] ^c[31] ^c[29] ^c[28] ^c[25] ^c[24] ^c[22] ^c[20] ^c[19] ^c[16] ^c[15] ^c[13] ^c[11] ^c[10] ^c[ 2] ^c[ 0] ;
            next_c[ 1] = d[ 1] ^c[30] ^c[26] ^c[25] ^c[24] ^c[21] ^c[17] ^c[16] ^c[15] ^c[12] ^c[ 8] ^c[ 7] ^c[ 5] ^c[ 4] ^c[ 2] ;
            next_c[ 0] = d[ 0] ^c[29] ^c[28] ^c[27] ^c[26] ^c[24] ^c[20] ^c[19] ^c[18] ^c[17] ^c[15] ^c[11] ^c[10] ^c[ 9] ^c[ 8] ^c[ 6] ^c[ 5] ^c[ 3] ^c[ 2] ;
            next_crc_140 = next_c;
        end
    endfunction

endmodule
