
module ecc_111_top

#

(

    parameter DATA_WIDTH = 111,

    parameter PARITY_WIDTH = 8

)

(

    input   [  DATA_WIDTH-1:0]   data_in,

    output  [  DATA_WIDTH-1:0]   data_out,

    input   [   PARITY_WIDTH-1:0]   parity_in,

    output  [   PARITY_WIDTH-1:0]   parity_out,

    input   bypass,

    output  reg [  DATA_WIDTH-1:0]   mask,

    output  sbit_err,

    output  dbit_err

);



wire  [   PARITY_WIDTH-1:0]   syndrome;

reg   [   1:0]              error;



assign parity_out = ecc_encode(data_in);

assign syndrome = parity_in ^ parity_out;

assign data_out = bypass ? data_in : data_in ^ mask;

assign sbit_err = bypass ? 1'b0 : error[0];

assign dbit_err = bypass ? 1'b0 : error[1];





always @(*)

begin

    error = 2'b00;

    case(syndrome)

    8'b00000000 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b00; end

    8'b10000011 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; error = 2'b01; end

    8'b10000101 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; error = 2'b01; end

    8'b10000110 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; error = 2'b01; end

    8'b00000111 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; error = 2'b01; end

    8'b10001001 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; error = 2'b01; end

    8'b10001010 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; error = 2'b01; end

    8'b00001011 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; error = 2'b01; end

    8'b10001100 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; error = 2'b01; end

    8'b00001101 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; error = 2'b01; end

    8'b00001110 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; error = 2'b01; end

    8'b10001111 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; error = 2'b01; end

    8'b10010001 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; error = 2'b01; end

    8'b10010010 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; error = 2'b01; end

    8'b00010011 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; error = 2'b01; end

    8'b10010100 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; error = 2'b01; end

    8'b00010101 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; error = 2'b01; end

    8'b00010110 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; error = 2'b01; end

    8'b10010111 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; error = 2'b01; end

    8'b10011000 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; error = 2'b01; end

    8'b00011001 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; error = 2'b01; end

    8'b00011010 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; error = 2'b01; end

    8'b10011011 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; error = 2'b01; end

    8'b00011100 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; error = 2'b01; end

    8'b10011101 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; error = 2'b01; end

    8'b10011110 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; error = 2'b01; end

    8'b00011111 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; error = 2'b01; end

    8'b10100001 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; error = 2'b01; end

    8'b10100010 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; error = 2'b01; end

    8'b00100011 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; error = 2'b01; end

    8'b10100100 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; error = 2'b01; end

    8'b00100101 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; error = 2'b01; end

    8'b00100110 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; error = 2'b01; end

    8'b10100111 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; error = 2'b01; end

    8'b10101000 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; error = 2'b01; end

    8'b00101001 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; error = 2'b01; end

    8'b00101010 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; error = 2'b01; end

    8'b10101011 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; error = 2'b01; end

    8'b00101100 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; error = 2'b01; end

    8'b10101101 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; error = 2'b01; end

    8'b10101110 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; error = 2'b01; end

    8'b00101111 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; error = 2'b01; end

    8'b10110000 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; error = 2'b01; end

    8'b00110001 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; error = 2'b01; end

    8'b00110010 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; error = 2'b01; end

    8'b10110011 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; error = 2'b01; end

    8'b00110100 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b10110101 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b10110110 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b00110111 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b00111000 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b10111001 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b10111010 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b00111011 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b10111100 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b00111101 : begin mask = 111'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b00111110 : begin mask = 111'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b10111111 : begin mask = 111'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11000001 : begin mask = 111'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11000010 : begin mask = 111'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01000011 : begin mask = 111'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11000100 : begin mask = 111'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01000101 : begin mask = 111'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01000110 : begin mask = 111'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11000111 : begin mask = 111'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11001000 : begin mask = 111'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01001001 : begin mask = 111'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01001010 : begin mask = 111'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11001011 : begin mask = 111'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01001100 : begin mask = 111'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11001101 : begin mask = 111'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11001110 : begin mask = 111'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01001111 : begin mask = 111'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11010000 : begin mask = 111'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01010001 : begin mask = 111'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01010010 : begin mask = 111'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11010011 : begin mask = 111'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01010100 : begin mask = 111'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11010101 : begin mask = 111'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11010110 : begin mask = 111'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01010111 : begin mask = 111'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01011000 : begin mask = 111'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11011001 : begin mask = 111'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11011010 : begin mask = 111'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01011011 : begin mask = 111'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11011100 : begin mask = 111'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01011101 : begin mask = 111'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01011110 : begin mask = 111'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11011111 : begin mask = 111'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11100000 : begin mask = 111'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01100001 : begin mask = 111'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01100010 : begin mask = 111'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11100011 : begin mask = 111'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01100100 : begin mask = 111'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11100101 : begin mask = 111'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11100110 : begin mask = 111'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01100111 : begin mask = 111'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01101000 : begin mask = 111'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11101001 : begin mask = 111'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11101010 : begin mask = 111'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01101011 : begin mask = 111'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11101100 : begin mask = 111'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01101101 : begin mask = 111'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01101110 : begin mask = 111'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11101111 : begin mask = 111'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01110000 : begin mask = 111'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11110001 : begin mask = 111'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11110010 : begin mask = 111'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01110011 : begin mask = 111'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b11110100 : begin mask = 111'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01110101 : begin mask = 111'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01110110 : begin mask = 111'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b10000000 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b01000000 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b00100000 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b00010000 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b00001000 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b00000100 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b00000010 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    8'b00000001 : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    default : begin mask = 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b10; end

    endcase

end



function [  PARITY_WIDTH-1:0] ecc_encode;

    input [ DATA_WIDTH-1:0] d;

    reg [ PARITY_WIDTH-1:0] p;

    begin

    p[0] = d[0] + d[1] + d[3] + d[4] + d[6] + d[8] + d[10] + d[11] + d[13] + d[15] + d[17] + d[19] + d[21] + d[23] + d[25] + d[26] + d[28] + d[30] + d[32] + d[34] + d[36] + d[38] + d[40] + d[42] + d[44] + d[46] + d[48] + d[50] + d[52] + d[54] + d[56] + d[57] + d[59] + d[61] + d[63] + d[65] + d[67] + d[69] + d[71] + d[73] + d[75] + d[77] + d[79] + d[81] + d[83] + d[85] + d[87] + d[89] + d[91] + d[93] + d[95] + d[97] + d[99] + d[101] + d[103] + d[105] + d[107] + d[109] ;

    p[1] = d[0] + d[2] + d[3] + d[5] + d[6] + d[9] + d[10] + d[12] + d[13] + d[16] + d[17] + d[20] + d[21] + d[24] + d[25] + d[27] + d[28] + d[31] + d[32] + d[35] + d[36] + d[39] + d[40] + d[43] + d[44] + d[47] + d[48] + d[51] + d[52] + d[55] + d[56] + d[58] + d[59] + d[62] + d[63] + d[66] + d[67] + d[70] + d[71] + d[74] + d[75] + d[78] + d[79] + d[82] + d[83] + d[86] + d[87] + d[90] + d[91] + d[94] + d[95] + d[98] + d[99] + d[102] + d[103] + d[106] + d[107] + d[110] ;

    p[2] = d[1] + d[2] + d[3] + d[7] + d[8] + d[9] + d[10] + d[14] + d[15] + d[16] + d[17] + d[22] + d[23] + d[24] + d[25] + d[29] + d[30] + d[31] + d[32] + d[37] + d[38] + d[39] + d[40] + d[45] + d[46] + d[47] + d[48] + d[53] + d[54] + d[55] + d[56] + d[60] + d[61] + d[62] + d[63] + d[68] + d[69] + d[70] + d[71] + d[76] + d[77] + d[78] + d[79] + d[84] + d[85] + d[86] + d[87] + d[92] + d[93] + d[94] + d[95] + d[100] + d[101] + d[102] + d[103] + d[108] + d[109] + d[110] ;

    p[3] = d[4] + d[5] + d[6] + d[7] + d[8] + d[9] + d[10] + d[18] + d[19] + d[20] + d[21] + d[22] + d[23] + d[24] + d[25] + d[33] + d[34] + d[35] + d[36] + d[37] + d[38] + d[39] + d[40] + d[49] + d[50] + d[51] + d[52] + d[53] + d[54] + d[55] + d[56] + d[64] + d[65] + d[66] + d[67] + d[68] + d[69] + d[70] + d[71] + d[80] + d[81] + d[82] + d[83] + d[84] + d[85] + d[86] + d[87] + d[96] + d[97] + d[98] + d[99] + d[100] + d[101] + d[102] + d[103] ;

    p[4] = d[11] + d[12] + d[13] + d[14] + d[15] + d[16] + d[17] + d[18] + d[19] + d[20] + d[21] + d[22] + d[23] + d[24] + d[25] + d[41] + d[42] + d[43] + d[44] + d[45] + d[46] + d[47] + d[48] + d[49] + d[50] + d[51] + d[52] + d[53] + d[54] + d[55] + d[56] + d[72] + d[73] + d[74] + d[75] + d[76] + d[77] + d[78] + d[79] + d[80] + d[81] + d[82] + d[83] + d[84] + d[85] + d[86] + d[87] + d[104] + d[105] + d[106] + d[107] + d[108] + d[109] + d[110] ;

    p[5] = d[26] + d[27] + d[28] + d[29] + d[30] + d[31] + d[32] + d[33] + d[34] + d[35] + d[36] + d[37] + d[38] + d[39] + d[40] + d[41] + d[42] + d[43] + d[44] + d[45] + d[46] + d[47] + d[48] + d[49] + d[50] + d[51] + d[52] + d[53] + d[54] + d[55] + d[56] + d[88] + d[89] + d[90] + d[91] + d[92] + d[93] + d[94] + d[95] + d[96] + d[97] + d[98] + d[99] + d[100] + d[101] + d[102] + d[103] + d[104] + d[105] + d[106] + d[107] + d[108] + d[109] + d[110] ;

    p[6] = d[57] + d[58] + d[59] + d[60] + d[61] + d[62] + d[63] + d[64] + d[65] + d[66] + d[67] + d[68] + d[69] + d[70] + d[71] + d[72] + d[73] + d[74] + d[75] + d[76] + d[77] + d[78] + d[79] + d[80] + d[81] + d[82] + d[83] + d[84] + d[85] + d[86] + d[87] + d[88] + d[89] + d[90] + d[91] + d[92] + d[93] + d[94] + d[95] + d[96] + d[97] + d[98] + d[99] + d[100] + d[101] + d[102] + d[103] + d[104] + d[105] + d[106] + d[107] + d[108] + d[109] + d[110] ;

    p[7] = d[0] + d[1] + d[2] + d[4] + d[5] + d[7] + d[10] + d[11] + d[12] + d[14] + d[17] + d[18] + d[21] + d[23] + d[24] + d[26] + d[27] + d[29] + d[32] + d[33] + d[36] + d[38] + d[39] + d[41] + d[44] + d[46] + d[47] + d[50] + d[51] + d[53] + d[56] + d[57] + d[58] + d[60] + d[63] + d[64] + d[67] + d[69] + d[70] + d[72] + d[75] + d[77] + d[78] + d[81] + d[82] + d[84] + d[87] + d[88] + d[91] + d[93] + d[94] + d[97] + d[98] + d[100] + d[103] + d[105] + d[106] + d[108] ;

    ecc_encode = p;

    end

endfunction



endmodule

