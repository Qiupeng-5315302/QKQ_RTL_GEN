
`timescale 1ns/1ps
module as6d_app_tb;

`include "APP_device_all_rtl_includes.vh"
`include "as6d_mep_all_includes.vh"
`include "wam_path_check_handle_app.sv"

    parameter   CSI2_DEVICE_VPG_BK_LINES_RS         = 10    ;    
    parameter   CSI2_DEVICE_VPG_DT_RS               =  6    ;
    parameter   CSI2_DEVICE_VPG_FRAME_NUM_MODE_RS   =  1    ;
    parameter   CSI2_DEVICE_VPG_HBP_TIME_RS         = 12    ;
    parameter   CSI2_DEVICE_VPG_HLINE_TIME_RS       = 15    ;
    parameter   CSI2_DEVICE_VPG_HSA_TIME_RS         = 12    ;
    parameter   CSI2_DEVICE_VPG_LINE_NUM_MODE_RS    =  2    ;
    parameter   CSI2_DEVICE_VPG_MAX_FRAME_NUM_RS    = 16    ;
    parameter   CSI2_DEVICE_VPG_PKT_SIZE_RS         = 14    ;
    parameter   CSI2_DEVICE_VPG_START_LINE_NUM_RS   = 16    ;
    parameter   CSI2_DEVICE_VPG_STEP_LINE_NUM_RS    = 16    ;
    parameter   CSI2_DEVICE_VPG_ACT_LINES_RS        = 14    ;
    parameter   CSI2_DEVICE_VPG_VBP_LINES_RS        = 10    ;
    parameter   CSI2_DEVICE_VPG_VC_RS               =  2    ;
    parameter   CSI2_DEVICE_VCX_DWIDTH              =  3    ;
    parameter   CSI2_DEVICE_VPG_VFP_LINES_RS        = 10    ;
    parameter   CSI2_DEVICE_VPG_VSA_LINES_RS        = 10    ;

`ifdef ASYNC_M1_4PIPE_CASE1
    `define ASYNC_M1
`elsif ASYNC_M1_8PIPE_CASE1
    `define ASYNC_M1
`elsif ASYNC_M1_8PIPE_CASE2
    `define ASYNC_M1
`elsif ASYNC_M2_2PIPE_CASE1
    `define ASYNC_M1
`elsif ASYNC_M2_4PIPE_CASE2
    `define ASYNC_M2
`endif

`ifdef DVP_RAW10_BYTELOC8
    `define DVP_RAW10
    `define AS6S_DVP
`elsif DVP_RAW10_BYTELOC7
    `define DVP_RAW10
    `define AS6S_DVP
`elsif DVP_RAW10_BYTELOC6
    `define DVP_RAW10
    `define AS6S_DVP
`elsif DVP_RAW10_BYTELOC5
    `define DVP_RAW10
    `define AS6S_DVP
`elsif DVP_RAW10_BYTELOC4
    `define DVP_RAW10
    `define AS6S_DVP
`elsif DVP_RAW10_BYTELOC3
    `define DVP_RAW10
    `define AS6S_DVP
`elsif DVP_RAW10_BYTELOC2
    `define DVP_RAW10
    `define AS6S_DVP
`elsif DVP_RAW10_BYTELOC1
    `define DVP_RAW10
    `define AS6S_DVP
`elsif DVP_RAW12_BYTELOC8
    `define DVP_RAW12
    `define AS6S_DVP
`elsif DVP_RAW12_BYTELOC7
    `define DVP_RAW12
    `define AS6S_DVP
`elsif DVP_RAW12_BYTELOC6
    `define DVP_RAW12
    `define AS6S_DVP
`elsif DVP_RAW12_BYTELOC5
    `define DVP_RAW12
    `define AS6S_DVP
`elsif DVP_RAW12_BYTELOC4
    `define DVP_RAW12
    `define AS6S_DVP
`elsif DVP_RAW12_BYTELOC3
    `define DVP_RAW12
    `define AS6S_DVP
`elsif DVP_RAW12_BYTELOC2
    `define DVP_RAW12
    `define AS6S_DVP
`elsif DVP_RAW12_BYTELOC1
    `define DVP_RAW12
    `define AS6S_DVP
`elsif DVP_RGB888_BYTELOC8
    `define DVP_RGB888
    `define AS6S_DVP
`elsif DVP_RGB888_BYTELOC7
    `define DVP_RGB888
    `define AS6S_DVP
`elsif DVP_RGB888_BYTELOC6
    `define DVP_RGB888
    `define AS6S_DVP
`elsif DVP_RGB888_BYTELOC5
    `define DVP_RGB888
    `define AS6S_DVP
`elsif DVP_RGB888_BYTELOC4
    `define DVP_RGB888
    `define AS6S_DVP
`elsif DVP_RGB888_BYTELOC3
    `define DVP_RGB888
    `define AS6S_DVP
`elsif DVP_RGB888_BYTELOC2
    `define DVP_RGB888
    `define AS6S_DVP
`elsif DVP_RGB888_BYTELOC1
    `define DVP_RGB888
    `define AS6S_DVP
`elsif DVP_YUV422_8BIT_UYVY
    `define DVP_YUV422_8BIT
    `define AS6S_DVP
`elsif DVP_YUV422_8BIT_YUYV
    `define DVP_YUV422_8BIT
    `define AS6S_DVP
`elsif DVP_YUV422_8BIT_YUYV_HS_TRIGGER
    `define DVP_YUV422_8BIT
    `define AS6S_DVP
`elsif DVP_RAW8
    `define AS6S_DVP
`elsif DVP_RGB565
    `define AS6S_DVP
`endif

wire clk_98M;
wire clk_99M;
wire clk_100M;
wire clk_101M;
wire clk_200M;
wire clk_1M;
wire clk_25M;
wire clk_10K;
wire clk_125M;

clk_generator#(100,1,1,"Mhz")clk_gen_100m(clk_100M);
clk_generator#(80 ,1,2,"Mhz")u0_clk_gen_100m(clk_98M);
clk_generator#(99 ,1,3,"Mhz")u1_clk_gen_100m(clk_99M);
clk_generator#(60,1,4,"Mhz")u3_clk_gen_100m(clk_101M);
clk_generator#(400,0,5,"Mhz")clk_gen_200m(clk_200M);
clk_generator#(1  ,0,6,"Mhz")clk_gen_1m(clk_1M);
clk_generator#(25,1,7,"Mhz")clk_gen_25m(clk_25M);
clk_generator#(10,1,8,"Khz")clk_gen_10k(clk_10K);
clk_generator#(125,1,9,"Mhz")clk_gen_125m(clk_125M);

reg                 clk_1M_rst_n;		// To u_as6d_app of as6d_app.v
reg                 reg_sync_aggr_0_video_mask_latch_reset;// To u_as6d_app of as6d_app.v
reg                 reg_sync_aggr_1_video_mask_latch_reset;// To u_as6d_app of as6d_app.v
reg                 reg_sync_aggr_2_video_mask_latch_reset;// To u_as6d_app of as6d_app.v
reg                 reg_sync_aggr_3_video_mask_latch_reset;// To u_as6d_app of as6d_app.v
reg [3:0]           reg_sync_aggr_auto_mask_en;// To u_as6d_app of as6d_app.v
reg                 reg_sync_aggr_check_framecount_en;// To u_as6d_app of as6d_app.v
reg                 reg_sync_aggr_check_linecount_en;// To u_as6d_app of as6d_app.v
reg [3:0]           reg_sync_aggr_force_video_mask;// To u_as6d_app of as6d_app.v
reg [3:0]           reg_sync_aggr_video_mask_restart;// To u_as6d_app of as6d_app.v
reg [5:0]           reg_sync_aggr_video_status_info_datatype;// To u_as6d_app of as6d_app.v
reg [15:0]          reg_sync_aggr_video_status_info_linecount;// To u_as6d_app of as6d_app.v
reg [4:0]           reg_sync_aggr_video_status_info_vc;// To u_as6d_app of as6d_app.v
reg [15:0]          reg_sync_aggr_video_status_info_wordcount;// To u_as6d_app of as6d_app.v
reg [19:0]          reg_sync_aggr_video_timeout_threshold;// To u_as6d_app of as6d_app.v

reg                 dvp_clk;        
reg                 dvp_clk_rst_n;        
reg                 test_mode;
reg    [6:0]        reg_mem_dt1_selz;
reg    [6:0]        reg_mem_dt2_selz;
reg    [6:0]        reg_mem_dt7_selz;
reg    [6:0]        reg_mem_dt8_selz;
reg    [7:0]        reg_mem_dt3_selz;
reg    [7:0]        reg_mem_dt4_selz;
reg                 reg_mem_dt3_selz_en;
reg                 reg_mem_dt4_selz_en;
reg    [7:0]        reg_vc_selz_l; 
reg    [7:0]        reg_vc_selz_h; 
reg                 treed_reg_bank_clk;
reg                 treed_reg_bank_clk_reset_n;
reg                 aggre_clk0;        
reg                 aggre_clk1;        
reg                 aggre_clk2;        
reg                 aggre_clk3;        
reg                 aggre_clk_rst_n0;    
reg                 aggre_clk_rst_n1;    
reg                 aggre_clk_rst_n2;    
reg                 aggre_clk_rst_n3;    
reg [15:0]          reg_app_sch0;        
reg [15:0]          reg_app_sch1;        
reg [15:0]          reg_app_sch2;        
reg [15:0]          reg_app_sch3;        
reg                 reg_sch0_frame_sync_lock;
reg                 reg_sch1_frame_sync_lock;
reg                 reg_sch2_frame_sync_lock;
reg                 reg_sch3_frame_sync_lock;
reg                 gpio2app_sch0_frame_sync_lock;
reg                 gpio2app_sch1_frame_sync_lock;
reg                 gpio2app_sch2_frame_sync_lock;
reg                 gpio2app_sch3_frame_sync_lock;
reg                 reg_app_sch0_frame_sync_lock;
reg                 reg_app_sch0_frame_sync_lock_force;
reg                 reg_app_sch1_frame_sync_lock;
reg                 reg_app_sch1_frame_sync_lock_force;
reg                 reg_app_sch2_frame_sync_lock;
reg                 reg_app_sch2_frame_sync_lock_force;
reg                 reg_app_sch3_frame_sync_lock;
reg                 reg_app_sch3_frame_sync_lock_force;

reg  [7:0]          reg_rd_pipe_fifo_full;
reg                 reg_all_pipe_wr_mode_strobe;
reg                 reg_app_aggregation_bypass;
reg                 reg_video_fifo_empty_depend_cnt_mux;
reg                 reg_delete_lp_depend_on_wc_mux;
reg                 reg_last_byte_header_down_mux; 
reg  [2:0]          reg_app_aggr0_vc_bit_override_en;
reg  [2:0]          reg_app_aggr0_vc_bit_override_value;
reg  [2:0]          reg_app_aggr1_vc_bit_override_en;
reg  [2:0]          reg_app_aggr1_vc_bit_override_value;
reg  [2:0]          reg_app_aggr2_vc_bit_override_en;
reg  [2:0]          reg_app_aggr2_vc_bit_override_value;
reg  [2:0]          reg_app_aggr3_vc_bit_override_en;
reg  [2:0]          reg_app_aggr3_vc_bit_override_value;
reg                 reg_app_vc_turn_over_en;
reg 	            reg_app_vc_turn_over_mode;

reg  [3:0]          reg_pipe_fifo_full_clear;
reg  [3:0]          reg_pipe_fifo_full_clear_last_four;
reg                 fifo_wrclk0;
reg                 fifo_rdclk0;
reg                 fifo_wrclk_rst_n0;
reg                 fifo_rdclk_rst_n0;
reg                 reg_line_delay_en0;
reg [1:0]           reg_pipe0_stream_sel;
reg [16:0]          reg_time_window0;
reg                 reg_video_loss_en0;
reg  [15:0]         reg_pipe0_map_en;            
reg  [3:0]          reg_pipe0_map0_aggr_id;            
reg  [3:0]          reg_pipe0_map1_aggr_id;            
reg  [3:0]          reg_pipe0_map2_aggr_id;            
reg  [3:0]          reg_pipe0_map3_aggr_id;            
reg  [3:0]          reg_pipe0_map4_aggr_id;            
reg  [3:0]          reg_pipe0_map5_aggr_id;            
reg  [3:0]          reg_pipe0_map6_aggr_id;            
reg  [3:0]          reg_pipe0_map7_aggr_id;            
reg  [3:0]          reg_pipe0_map8_aggr_id;            
reg  [3:0]          reg_pipe0_map9_aggr_id;            
reg  [3:0]          reg_pipe0_map10_aggr_id;            
reg  [3:0]          reg_pipe0_map11_aggr_id;            
reg  [3:0]          reg_pipe0_map12_aggr_id;            
reg  [3:0]          reg_pipe0_map13_aggr_id;            
reg  [3:0]          reg_pipe0_map14_aggr_id;            
reg  [3:0]          reg_pipe0_map15_aggr_id;            
reg  [1:0]          reg_pipe0_map0_vc_source;            
reg  [1:0]          reg_pipe0_map1_vc_source;            
reg  [1:0]          reg_pipe0_map2_vc_source;            
reg  [1:0]          reg_pipe0_map3_vc_source;            
reg  [1:0]          reg_pipe0_map4_vc_source;            
reg  [1:0]          reg_pipe0_map5_vc_source;            
reg  [1:0]          reg_pipe0_map6_vc_source;            
reg  [1:0]          reg_pipe0_map7_vc_source;            
reg  [1:0]          reg_pipe0_map8_vc_source;            
reg  [1:0]          reg_pipe0_map9_vc_source;            
reg  [1:0]          reg_pipe0_map10_vc_source;            
reg  [1:0]          reg_pipe0_map11_vc_source;            
reg  [1:0]          reg_pipe0_map12_vc_source;            
reg  [1:0]          reg_pipe0_map13_vc_source;            
reg  [1:0]          reg_pipe0_map14_vc_source;            
reg  [1:0]          reg_pipe0_map15_vc_source;            
reg  [1:0]          reg_pipe0_map0_vc_dest;            
reg  [1:0]          reg_pipe0_map1_vc_dest;            
reg  [1:0]          reg_pipe0_map2_vc_dest;            
reg  [1:0]          reg_pipe0_map3_vc_dest;            
reg  [1:0]          reg_pipe0_map4_vc_dest;            
reg  [1:0]          reg_pipe0_map5_vc_dest;            
reg  [1:0]          reg_pipe0_map6_vc_dest;            
reg  [1:0]          reg_pipe0_map7_vc_dest;            
reg  [1:0]          reg_pipe0_map8_vc_dest;            
reg  [1:0]          reg_pipe0_map9_vc_dest;            
reg  [1:0]          reg_pipe0_map10_vc_dest;            
reg  [1:0]          reg_pipe0_map11_vc_dest;            
reg  [1:0]          reg_pipe0_map12_vc_dest;            
reg  [1:0]          reg_pipe0_map13_vc_dest;            
reg  [1:0]          reg_pipe0_map14_vc_dest;            
reg  [1:0]          reg_pipe0_map15_vc_dest;            
reg  [5:0]          reg_pipe0_map0_dt_source;            
reg  [5:0]          reg_pipe0_map1_dt_source;            
reg  [5:0]          reg_pipe0_map2_dt_source;            
reg  [5:0]          reg_pipe0_map3_dt_source;            
reg  [5:0]          reg_pipe0_map4_dt_source;            
reg  [5:0]          reg_pipe0_map5_dt_source;            
reg  [5:0]          reg_pipe0_map6_dt_source;            
reg  [5:0]          reg_pipe0_map7_dt_source;            
reg  [5:0]          reg_pipe0_map8_dt_source;            
reg  [5:0]          reg_pipe0_map9_dt_source;            
reg  [5:0]          reg_pipe0_map10_dt_source;            
reg  [5:0]          reg_pipe0_map11_dt_source;            
reg  [5:0]          reg_pipe0_map12_dt_source;            
reg  [5:0]          reg_pipe0_map13_dt_source;            
reg  [5:0]          reg_pipe0_map14_dt_source;            
reg  [5:0]          reg_pipe0_map15_dt_source;            
reg  [5:0]          reg_pipe0_map0_dt_dest;            
reg  [5:0]          reg_pipe0_map1_dt_dest;            
reg  [5:0]          reg_pipe0_map2_dt_dest;            
reg  [5:0]          reg_pipe0_map3_dt_dest;            
reg  [5:0]          reg_pipe0_map4_dt_dest;            
reg  [5:0]          reg_pipe0_map5_dt_dest;            
reg  [5:0]          reg_pipe0_map6_dt_dest;            
reg  [5:0]          reg_pipe0_map7_dt_dest;            
reg  [5:0]          reg_pipe0_map8_dt_dest;            
reg  [5:0]          reg_pipe0_map9_dt_dest;            
reg  [5:0]          reg_pipe0_map10_dt_dest;            
reg  [5:0]          reg_pipe0_map11_dt_dest;            
reg  [5:0]          reg_pipe0_map12_dt_dest;            
reg  [5:0]          reg_pipe0_map13_dt_dest;            
reg  [5:0]          reg_pipe0_map14_dt_dest;            
reg  [5:0]          reg_pipe0_map15_dt_dest;            
reg  [1:0]          reg_pipe0_wr_mode;
wire [31:0]         reg_rd_app_full_cnt_async_fifo_pipe0;
wire [31:0]         reg_rd_app_full_cnt_sync_fifo_pipe0;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_pf_pipe0;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_ph_pipe0;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fe_pipe0;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fs_pipe0;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_le_pipe0;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_ls_pipe0;
reg                 reg_clear_app_full_cnt_async_fifo_pipe0;
reg                 reg_clear_app_full_cnt_sync_fifo_pipe0;
reg                 reg_clear_resv_pkt_cnt_lp_pf_pipe0;
reg                 reg_clear_resv_pkt_cnt_lp_ph_pipe0;
reg                 reg_clear_resv_pkt_cnt_sp_fe_pipe0;
reg                 reg_clear_resv_pkt_cnt_sp_fs_pipe0;
reg                 reg_clear_resv_pkt_cnt_sp_le_pipe0;
reg                 reg_clear_resv_pkt_cnt_sp_ls_pipe0;
reg                 fifo_wrclk1;
reg                 fifo_rdclk1;
reg                 fifo_wrclk_rst_n1;
reg                 fifo_rdclk_rst_n1;
reg                 reg_line_delay_en1;
reg [1:0]           reg_pipe1_stream_sel;
reg [16:0]          reg_time_window1;
reg                 reg_video_loss_en1;
reg  [15:0]         reg_pipe1_map_en;            
reg  [3:0]          reg_pipe1_map0_aggr_id;            
reg  [3:0]          reg_pipe1_map1_aggr_id;            
reg  [3:0]          reg_pipe1_map2_aggr_id;            
reg  [3:0]          reg_pipe1_map3_aggr_id;            
reg  [3:0]          reg_pipe1_map4_aggr_id;            
reg  [3:0]          reg_pipe1_map5_aggr_id;            
reg  [3:0]          reg_pipe1_map6_aggr_id;            
reg  [3:0]          reg_pipe1_map7_aggr_id;            
reg  [3:0]          reg_pipe1_map8_aggr_id;            
reg  [3:0]          reg_pipe1_map9_aggr_id;            
reg  [3:0]          reg_pipe1_map10_aggr_id;            
reg  [3:0]          reg_pipe1_map11_aggr_id;            
reg  [3:0]          reg_pipe1_map12_aggr_id;            
reg  [3:0]          reg_pipe1_map13_aggr_id;            
reg  [3:0]          reg_pipe1_map14_aggr_id;            
reg  [3:0]          reg_pipe1_map15_aggr_id;            
reg  [1:0]          reg_pipe1_map0_vc_source;            
reg  [1:0]          reg_pipe1_map1_vc_source;            
reg  [1:0]          reg_pipe1_map2_vc_source;            
reg  [1:0]          reg_pipe1_map3_vc_source;            
reg  [1:0]          reg_pipe1_map4_vc_source;            
reg  [1:0]          reg_pipe1_map5_vc_source;            
reg  [1:0]          reg_pipe1_map6_vc_source;            
reg  [1:0]          reg_pipe1_map7_vc_source;            
reg  [1:0]          reg_pipe1_map8_vc_source;            
reg  [1:0]          reg_pipe1_map9_vc_source;            
reg  [1:0]          reg_pipe1_map10_vc_source;            
reg  [1:0]          reg_pipe1_map11_vc_source;            
reg  [1:0]          reg_pipe1_map12_vc_source;            
reg  [1:0]          reg_pipe1_map13_vc_source;            
reg  [1:0]          reg_pipe1_map14_vc_source;            
reg  [1:0]          reg_pipe1_map15_vc_source;            
reg  [1:0]          reg_pipe1_map0_vc_dest;            
reg  [1:0]          reg_pipe1_map1_vc_dest;            
reg  [1:0]          reg_pipe1_map2_vc_dest;            
reg  [1:0]          reg_pipe1_map3_vc_dest;            
reg  [1:0]          reg_pipe1_map4_vc_dest;            
reg  [1:0]          reg_pipe1_map5_vc_dest;            
reg  [1:0]          reg_pipe1_map6_vc_dest;            
reg  [1:0]          reg_pipe1_map7_vc_dest;            
reg  [1:0]          reg_pipe1_map8_vc_dest;            
reg  [1:0]          reg_pipe1_map9_vc_dest;            
reg  [1:0]          reg_pipe1_map10_vc_dest;            
reg  [1:0]          reg_pipe1_map11_vc_dest;            
reg  [1:0]          reg_pipe1_map12_vc_dest;            
reg  [1:0]          reg_pipe1_map13_vc_dest;            
reg  [1:0]          reg_pipe1_map14_vc_dest;            
reg  [1:0]          reg_pipe1_map15_vc_dest;            
reg  [5:0]          reg_pipe1_map0_dt_source;            
reg  [5:0]          reg_pipe1_map1_dt_source;            
reg  [5:0]          reg_pipe1_map2_dt_source;            
reg  [5:0]          reg_pipe1_map3_dt_source;            
reg  [5:0]          reg_pipe1_map4_dt_source;            
reg  [5:0]          reg_pipe1_map5_dt_source;            
reg  [5:0]          reg_pipe1_map6_dt_source;            
reg  [5:0]          reg_pipe1_map7_dt_source;            
reg  [5:0]          reg_pipe1_map8_dt_source;            
reg  [5:0]          reg_pipe1_map9_dt_source;            
reg  [5:0]          reg_pipe1_map10_dt_source;            
reg  [5:0]          reg_pipe1_map11_dt_source;            
reg  [5:0]          reg_pipe1_map12_dt_source;            
reg  [5:0]          reg_pipe1_map13_dt_source;            
reg  [5:0]          reg_pipe1_map14_dt_source;            
reg  [5:0]          reg_pipe1_map15_dt_source;            
reg  [5:0]          reg_pipe1_map0_dt_dest;            
reg  [5:0]          reg_pipe1_map1_dt_dest;            
reg  [5:0]          reg_pipe1_map2_dt_dest;            
reg  [5:0]          reg_pipe1_map3_dt_dest;            
reg  [5:0]          reg_pipe1_map4_dt_dest;            
reg  [5:0]          reg_pipe1_map5_dt_dest;            
reg  [5:0]          reg_pipe1_map6_dt_dest;            
reg  [5:0]          reg_pipe1_map7_dt_dest;            
reg  [5:0]          reg_pipe1_map8_dt_dest;            
reg  [5:0]          reg_pipe1_map9_dt_dest;            
reg  [5:0]          reg_pipe1_map10_dt_dest;            
reg  [5:0]          reg_pipe1_map11_dt_dest;            
reg  [5:0]          reg_pipe1_map12_dt_dest;            
reg  [5:0]          reg_pipe1_map13_dt_dest;            
reg  [5:0]          reg_pipe1_map14_dt_dest;            
reg  [5:0]          reg_pipe1_map15_dt_dest;            
reg  [1:0]          reg_pipe1_wr_mode;
wire [31:0]         reg_rd_app_full_cnt_async_fifo_pipe1;
wire [31:0]         reg_rd_app_full_cnt_sync_fifo_pipe1;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_pf_pipe1;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_ph_pipe1;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fe_pipe1;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fs_pipe1;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_le_pipe1;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_ls_pipe1;
reg                 reg_clear_app_full_cnt_async_fifo_pipe1;
reg                 reg_clear_app_full_cnt_sync_fifo_pipe1;
reg                 reg_clear_resv_pkt_cnt_lp_pf_pipe1 ;
reg                 reg_clear_resv_pkt_cnt_lp_ph_pipe1 ;
reg                 reg_clear_resv_pkt_cnt_sp_fe_pipe1 ;
reg                 reg_clear_resv_pkt_cnt_sp_fs_pipe1 ;
reg                 reg_clear_resv_pkt_cnt_sp_le_pipe1 ;
reg                 reg_clear_resv_pkt_cnt_sp_ls_pipe1 ;
reg                 fifo_wrclk2;
reg                 fifo_rdclk2;
reg                 fifo_wrclk_rst_n2;
reg                 fifo_rdclk_rst_n2;
reg                 reg_line_delay_en2;
reg [1:0]           reg_pipe2_stream_sel;
reg [16:0]          reg_time_window2;
reg                 reg_video_loss_en2;
reg  [15:0]         reg_pipe2_map_en;            
reg  [3:0]          reg_pipe2_map0_aggr_id;            
reg  [3:0]          reg_pipe2_map1_aggr_id;            
reg  [3:0]          reg_pipe2_map2_aggr_id;            
reg  [3:0]          reg_pipe2_map3_aggr_id;            
reg  [3:0]          reg_pipe2_map4_aggr_id;            
reg  [3:0]          reg_pipe2_map5_aggr_id;            
reg  [3:0]          reg_pipe2_map6_aggr_id;            
reg  [3:0]          reg_pipe2_map7_aggr_id;            
reg  [3:0]          reg_pipe2_map8_aggr_id;            
reg  [3:0]          reg_pipe2_map9_aggr_id;            
reg  [3:0]          reg_pipe2_map10_aggr_id;            
reg  [3:0]          reg_pipe2_map11_aggr_id;            
reg  [3:0]          reg_pipe2_map12_aggr_id;            
reg  [3:0]          reg_pipe2_map13_aggr_id;            
reg  [3:0]          reg_pipe2_map14_aggr_id;            
reg  [3:0]          reg_pipe2_map15_aggr_id;            
reg  [1:0]          reg_pipe2_map0_vc_source;            
reg  [1:0]          reg_pipe2_map1_vc_source;            
reg  [1:0]          reg_pipe2_map2_vc_source;            
reg  [1:0]          reg_pipe2_map3_vc_source;            
reg  [1:0]          reg_pipe2_map4_vc_source;            
reg  [1:0]          reg_pipe2_map5_vc_source;            
reg  [1:0]          reg_pipe2_map6_vc_source;            
reg  [1:0]          reg_pipe2_map7_vc_source;            
reg  [1:0]          reg_pipe2_map8_vc_source;            
reg  [1:0]          reg_pipe2_map9_vc_source;            
reg  [1:0]          reg_pipe2_map10_vc_source;            
reg  [1:0]          reg_pipe2_map11_vc_source;            
reg  [1:0]          reg_pipe2_map12_vc_source;            
reg  [1:0]          reg_pipe2_map13_vc_source;            
reg  [1:0]          reg_pipe2_map14_vc_source;            
reg  [1:0]          reg_pipe2_map15_vc_source;            
reg  [1:0]          reg_pipe2_map0_vc_dest;            
reg  [1:0]          reg_pipe2_map1_vc_dest;            
reg  [1:0]          reg_pipe2_map2_vc_dest;            
reg  [1:0]          reg_pipe2_map3_vc_dest;            
reg  [1:0]          reg_pipe2_map4_vc_dest;            
reg  [1:0]          reg_pipe2_map5_vc_dest;            
reg  [1:0]          reg_pipe2_map6_vc_dest;            
reg  [1:0]          reg_pipe2_map7_vc_dest;            
reg  [1:0]          reg_pipe2_map8_vc_dest;            
reg  [1:0]          reg_pipe2_map9_vc_dest;            
reg  [1:0]          reg_pipe2_map10_vc_dest;            
reg  [1:0]          reg_pipe2_map11_vc_dest;            
reg  [1:0]          reg_pipe2_map12_vc_dest;            
reg  [1:0]          reg_pipe2_map13_vc_dest;            
reg  [1:0]          reg_pipe2_map14_vc_dest;            
reg  [1:0]          reg_pipe2_map15_vc_dest;            
reg  [5:0]          reg_pipe2_map0_dt_source;            
reg  [5:0]          reg_pipe2_map1_dt_source;            
reg  [5:0]          reg_pipe2_map2_dt_source;            
reg  [5:0]          reg_pipe2_map3_dt_source;            
reg  [5:0]          reg_pipe2_map4_dt_source;            
reg  [5:0]          reg_pipe2_map5_dt_source;            
reg  [5:0]          reg_pipe2_map6_dt_source;            
reg  [5:0]          reg_pipe2_map7_dt_source;            
reg  [5:0]          reg_pipe2_map8_dt_source;            
reg  [5:0]          reg_pipe2_map9_dt_source;            
reg  [5:0]          reg_pipe2_map10_dt_source;            
reg  [5:0]          reg_pipe2_map11_dt_source;            
reg  [5:0]          reg_pipe2_map12_dt_source;            
reg  [5:0]          reg_pipe2_map13_dt_source;            
reg  [5:0]          reg_pipe2_map14_dt_source;            
reg  [5:0]          reg_pipe2_map15_dt_source;            
reg  [5:0]          reg_pipe2_map0_dt_dest;            
reg  [5:0]          reg_pipe2_map1_dt_dest;            
reg  [5:0]          reg_pipe2_map2_dt_dest;            
reg  [5:0]          reg_pipe2_map3_dt_dest;            
reg  [5:0]          reg_pipe2_map4_dt_dest;            
reg  [5:0]          reg_pipe2_map5_dt_dest;            
reg  [5:0]          reg_pipe2_map6_dt_dest;            
reg  [5:0]          reg_pipe2_map7_dt_dest;            
reg  [5:0]          reg_pipe2_map8_dt_dest;            
reg  [5:0]          reg_pipe2_map9_dt_dest;            
reg  [5:0]          reg_pipe2_map10_dt_dest;            
reg  [5:0]          reg_pipe2_map11_dt_dest;            
reg  [5:0]          reg_pipe2_map12_dt_dest;            
reg  [5:0]          reg_pipe2_map13_dt_dest;            
reg  [5:0]          reg_pipe2_map14_dt_dest;            
reg  [5:0]          reg_pipe2_map15_dt_dest;            
reg  [1:0]          reg_pipe2_wr_mode;
wire [31:0]         reg_rd_app_full_cnt_async_fifo_pipe2;
wire [31:0]         reg_rd_app_full_cnt_sync_fifo_pipe2;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_pf_pipe2;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_ph_pipe2;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fe_pipe2;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fs_pipe2;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_le_pipe2;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_ls_pipe2;
reg                reg_clear_app_full_cnt_async_fifo_pipe2;
reg                reg_clear_app_full_cnt_sync_fifo_pipe2;
reg                reg_clear_resv_pkt_cnt_lp_pf_pipe2 ;
reg                reg_clear_resv_pkt_cnt_lp_ph_pipe2 ;
reg                reg_clear_resv_pkt_cnt_sp_fe_pipe2 ;
reg                reg_clear_resv_pkt_cnt_sp_fs_pipe2 ;
reg                reg_clear_resv_pkt_cnt_sp_le_pipe2 ;
reg                reg_clear_resv_pkt_cnt_sp_ls_pipe2 ;
reg                 fifo_wrclk3;
reg                 fifo_rdclk3;
reg                 fifo_wrclk_rst_n3;
reg                 fifo_rdclk_rst_n3;
reg                 reg_line_delay_en3;
reg [1:0]           reg_pipe3_stream_sel;
reg [16:0]          reg_time_window3;
reg                 reg_video_loss_en3;
reg  [15:0]         reg_pipe3_map_en;            
reg  [3:0]          reg_pipe3_map0_aggr_id;            
reg  [3:0]          reg_pipe3_map1_aggr_id;            
reg  [3:0]          reg_pipe3_map2_aggr_id;            
reg  [3:0]          reg_pipe3_map3_aggr_id;            
reg  [3:0]          reg_pipe3_map4_aggr_id;            
reg  [3:0]          reg_pipe3_map5_aggr_id;            
reg  [3:0]          reg_pipe3_map6_aggr_id;            
reg  [3:0]          reg_pipe3_map7_aggr_id;            
reg  [3:0]          reg_pipe3_map8_aggr_id;            
reg  [3:0]          reg_pipe3_map9_aggr_id;            
reg  [3:0]          reg_pipe3_map10_aggr_id;            
reg  [3:0]          reg_pipe3_map11_aggr_id;            
reg  [3:0]          reg_pipe3_map12_aggr_id;            
reg  [3:0]          reg_pipe3_map13_aggr_id;            
reg  [3:0]          reg_pipe3_map14_aggr_id;            
reg  [3:0]          reg_pipe3_map15_aggr_id;            
reg  [1:0]          reg_pipe3_map0_vc_source;            
reg  [1:0]          reg_pipe3_map1_vc_source;            
reg  [1:0]          reg_pipe3_map2_vc_source;            
reg  [1:0]          reg_pipe3_map3_vc_source;            
reg  [1:0]          reg_pipe3_map4_vc_source;            
reg  [1:0]          reg_pipe3_map5_vc_source;            
reg  [1:0]          reg_pipe3_map6_vc_source;            
reg  [1:0]          reg_pipe3_map7_vc_source;            
reg  [1:0]          reg_pipe3_map8_vc_source;            
reg  [1:0]          reg_pipe3_map9_vc_source;            
reg  [1:0]          reg_pipe3_map10_vc_source;            
reg  [1:0]          reg_pipe3_map11_vc_source;            
reg  [1:0]          reg_pipe3_map12_vc_source;            
reg  [1:0]          reg_pipe3_map13_vc_source;            
reg  [1:0]          reg_pipe3_map14_vc_source;            
reg  [1:0]          reg_pipe3_map15_vc_source;            
reg  [1:0]          reg_pipe3_map0_vc_dest;            
reg  [1:0]          reg_pipe3_map1_vc_dest;            
reg  [1:0]          reg_pipe3_map2_vc_dest;            
reg  [1:0]          reg_pipe3_map3_vc_dest;            
reg  [1:0]          reg_pipe3_map4_vc_dest;            
reg  [1:0]          reg_pipe3_map5_vc_dest;            
reg  [1:0]          reg_pipe3_map6_vc_dest;            
reg  [1:0]          reg_pipe3_map7_vc_dest;            
reg  [1:0]          reg_pipe3_map8_vc_dest;            
reg  [1:0]          reg_pipe3_map9_vc_dest;            
reg  [1:0]          reg_pipe3_map10_vc_dest;            
reg  [1:0]          reg_pipe3_map11_vc_dest;            
reg  [1:0]          reg_pipe3_map12_vc_dest;            
reg  [1:0]          reg_pipe3_map13_vc_dest;            
reg  [1:0]          reg_pipe3_map14_vc_dest;            
reg  [1:0]          reg_pipe3_map15_vc_dest;            
reg  [5:0]          reg_pipe3_map0_dt_source;            
reg  [5:0]          reg_pipe3_map1_dt_source;            
reg  [5:0]          reg_pipe3_map2_dt_source;            
reg  [5:0]          reg_pipe3_map3_dt_source;            
reg  [5:0]          reg_pipe3_map4_dt_source;            
reg  [5:0]          reg_pipe3_map5_dt_source;            
reg  [5:0]          reg_pipe3_map6_dt_source;            
reg  [5:0]          reg_pipe3_map7_dt_source;            
reg  [5:0]          reg_pipe3_map8_dt_source;            
reg  [5:0]          reg_pipe3_map9_dt_source;            
reg  [5:0]          reg_pipe3_map10_dt_source;            
reg  [5:0]          reg_pipe3_map11_dt_source;            
reg  [5:0]          reg_pipe3_map12_dt_source;            
reg  [5:0]          reg_pipe3_map13_dt_source;            
reg  [5:0]          reg_pipe3_map14_dt_source;            
reg  [5:0]          reg_pipe3_map15_dt_source;            
reg  [5:0]          reg_pipe3_map0_dt_dest;            
reg  [5:0]          reg_pipe3_map1_dt_dest;            
reg  [5:0]          reg_pipe3_map2_dt_dest;            
reg  [5:0]          reg_pipe3_map3_dt_dest;            
reg  [5:0]          reg_pipe3_map4_dt_dest;            
reg  [5:0]          reg_pipe3_map5_dt_dest;            
reg  [5:0]          reg_pipe3_map6_dt_dest;            
reg  [5:0]          reg_pipe3_map7_dt_dest;            
reg  [5:0]          reg_pipe3_map8_dt_dest;            
reg  [5:0]          reg_pipe3_map9_dt_dest;            
reg  [5:0]          reg_pipe3_map10_dt_dest;            
reg  [5:0]          reg_pipe3_map11_dt_dest;            
reg  [5:0]          reg_pipe3_map12_dt_dest;            
reg  [5:0]          reg_pipe3_map13_dt_dest;            
reg  [5:0]          reg_pipe3_map14_dt_dest;            
reg  [5:0]          reg_pipe3_map15_dt_dest;            
reg  [1:0]          reg_pipe3_wr_mode;
wire [31:0]         reg_rd_app_full_cnt_async_fifo_pipe3;
wire [31:0]         reg_rd_app_full_cnt_sync_fifo_pipe3;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_pf_pipe3;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_ph_pipe3;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fe_pipe3;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fs_pipe3;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_le_pipe3;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_ls_pipe3;
reg                reg_clear_app_full_cnt_async_fifo_pipe3;
reg                reg_clear_app_full_cnt_sync_fifo_pipe3;
reg                reg_clear_resv_pkt_cnt_lp_pf_pipe3 ;
reg                reg_clear_resv_pkt_cnt_lp_ph_pipe3 ;
reg                reg_clear_resv_pkt_cnt_sp_fe_pipe3 ;
reg                reg_clear_resv_pkt_cnt_sp_fs_pipe3 ;
reg                reg_clear_resv_pkt_cnt_sp_le_pipe3 ;
reg                reg_clear_resv_pkt_cnt_sp_ls_pipe3 ;
reg                 fifo_wrclk4;
reg                 fifo_rdclk4;
reg                 fifo_wrclk_rst_n4;
reg                 fifo_rdclk_rst_n4;
reg                 reg_line_delay_en4;
reg [1:0]           reg_pipe4_stream_sel;
reg [16:0]          reg_time_window4;
reg                 reg_video_loss_en4;
reg  [15:0]         reg_pipe4_map_en;            
reg  [3:0]          reg_pipe4_map0_aggr_id;            
reg  [3:0]          reg_pipe4_map1_aggr_id;            
reg  [3:0]          reg_pipe4_map2_aggr_id;            
reg  [3:0]          reg_pipe4_map3_aggr_id;            
reg  [3:0]          reg_pipe4_map4_aggr_id;            
reg  [3:0]          reg_pipe4_map5_aggr_id;            
reg  [3:0]          reg_pipe4_map6_aggr_id;            
reg  [3:0]          reg_pipe4_map7_aggr_id;            
reg  [3:0]          reg_pipe4_map8_aggr_id;            
reg  [3:0]          reg_pipe4_map9_aggr_id;            
reg  [3:0]          reg_pipe4_map10_aggr_id;            
reg  [3:0]          reg_pipe4_map11_aggr_id;            
reg  [3:0]          reg_pipe4_map12_aggr_id;            
reg  [3:0]          reg_pipe4_map13_aggr_id;            
reg  [3:0]          reg_pipe4_map14_aggr_id;            
reg  [3:0]          reg_pipe4_map15_aggr_id;            
reg  [1:0]          reg_pipe4_map0_vc_source;            
reg  [1:0]          reg_pipe4_map1_vc_source;            
reg  [1:0]          reg_pipe4_map2_vc_source;            
reg  [1:0]          reg_pipe4_map3_vc_source;            
reg  [1:0]          reg_pipe4_map4_vc_source;            
reg  [1:0]          reg_pipe4_map5_vc_source;            
reg  [1:0]          reg_pipe4_map6_vc_source;            
reg  [1:0]          reg_pipe4_map7_vc_source;            
reg  [1:0]          reg_pipe4_map8_vc_source;            
reg  [1:0]          reg_pipe4_map9_vc_source;            
reg  [1:0]          reg_pipe4_map10_vc_source;            
reg  [1:0]          reg_pipe4_map11_vc_source;            
reg  [1:0]          reg_pipe4_map12_vc_source;            
reg  [1:0]          reg_pipe4_map13_vc_source;            
reg  [1:0]          reg_pipe4_map14_vc_source;            
reg  [1:0]          reg_pipe4_map15_vc_source;            
reg  [1:0]          reg_pipe4_map0_vc_dest;            
reg  [1:0]          reg_pipe4_map1_vc_dest;            
reg  [1:0]          reg_pipe4_map2_vc_dest;            
reg  [1:0]          reg_pipe4_map3_vc_dest;            
reg  [1:0]          reg_pipe4_map4_vc_dest;            
reg  [1:0]          reg_pipe4_map5_vc_dest;            
reg  [1:0]          reg_pipe4_map6_vc_dest;            
reg  [1:0]          reg_pipe4_map7_vc_dest;            
reg  [1:0]          reg_pipe4_map8_vc_dest;            
reg  [1:0]          reg_pipe4_map9_vc_dest;            
reg  [1:0]          reg_pipe4_map10_vc_dest;            
reg  [1:0]          reg_pipe4_map11_vc_dest;            
reg  [1:0]          reg_pipe4_map12_vc_dest;            
reg  [1:0]          reg_pipe4_map13_vc_dest;            
reg  [1:0]          reg_pipe4_map14_vc_dest;            
reg  [1:0]          reg_pipe4_map15_vc_dest;            
reg  [5:0]          reg_pipe4_map0_dt_source;            
reg  [5:0]          reg_pipe4_map1_dt_source;            
reg  [5:0]          reg_pipe4_map2_dt_source;            
reg  [5:0]          reg_pipe4_map3_dt_source;            
reg  [5:0]          reg_pipe4_map4_dt_source;            
reg  [5:0]          reg_pipe4_map5_dt_source;            
reg  [5:0]          reg_pipe4_map6_dt_source;            
reg  [5:0]          reg_pipe4_map7_dt_source;            
reg  [5:0]          reg_pipe4_map8_dt_source;            
reg  [5:0]          reg_pipe4_map9_dt_source;            
reg  [5:0]          reg_pipe4_map10_dt_source;            
reg  [5:0]          reg_pipe4_map11_dt_source;            
reg  [5:0]          reg_pipe4_map12_dt_source;            
reg  [5:0]          reg_pipe4_map13_dt_source;            
reg  [5:0]          reg_pipe4_map14_dt_source;            
reg  [5:0]          reg_pipe4_map15_dt_source;            
reg  [5:0]          reg_pipe4_map0_dt_dest;            
reg  [5:0]          reg_pipe4_map1_dt_dest;            
reg  [5:0]          reg_pipe4_map2_dt_dest;            
reg  [5:0]          reg_pipe4_map3_dt_dest;            
reg  [5:0]          reg_pipe4_map4_dt_dest;            
reg  [5:0]          reg_pipe4_map5_dt_dest;            
reg  [5:0]          reg_pipe4_map6_dt_dest;            
reg  [5:0]          reg_pipe4_map7_dt_dest;            
reg  [5:0]          reg_pipe4_map8_dt_dest;            
reg  [5:0]          reg_pipe4_map9_dt_dest;            
reg  [5:0]          reg_pipe4_map10_dt_dest;            
reg  [5:0]          reg_pipe4_map11_dt_dest;            
reg  [5:0]          reg_pipe4_map12_dt_dest;            
reg  [5:0]          reg_pipe4_map13_dt_dest;            
reg  [5:0]          reg_pipe4_map14_dt_dest;            
reg  [5:0]          reg_pipe4_map15_dt_dest;            
reg  [1:0]          reg_pipe4_wr_mode;
wire [31:0]         reg_rd_app_full_cnt_async_fifo_pipe4;
wire [31:0]         reg_rd_app_full_cnt_sync_fifo_pipe4;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_pf_pipe4;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_ph_pipe4;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fe_pipe4;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fs_pipe4;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_le_pipe4;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_ls_pipe4;
reg                reg_clear_app_full_cnt_async_fifo_pipe4;
reg                reg_clear_app_full_cnt_sync_fifo_pipe4;
reg                reg_clear_resv_pkt_cnt_lp_pf_pipe4 ;
reg                reg_clear_resv_pkt_cnt_lp_ph_pipe4 ;
reg                reg_clear_resv_pkt_cnt_sp_fe_pipe4 ;
reg                reg_clear_resv_pkt_cnt_sp_fs_pipe4 ;
reg                reg_clear_resv_pkt_cnt_sp_le_pipe4 ;
reg                reg_clear_resv_pkt_cnt_sp_ls_pipe4 ;
reg                 fifo_wrclk5;
reg                 fifo_rdclk5;
reg                 fifo_wrclk_rst_n5;
reg                 fifo_rdclk_rst_n5;
reg                 reg_line_delay_en5;
reg [1:0]           reg_pipe5_stream_sel;
reg [16:0]          reg_time_window5;
reg                 reg_video_loss_en5;
reg  [15:0]         reg_pipe5_map_en;            
reg  [3:0]          reg_pipe5_map0_aggr_id;            
reg  [3:0]          reg_pipe5_map1_aggr_id;            
reg  [3:0]          reg_pipe5_map2_aggr_id;            
reg  [3:0]          reg_pipe5_map3_aggr_id;            
reg  [3:0]          reg_pipe5_map4_aggr_id;            
reg  [3:0]          reg_pipe5_map5_aggr_id;            
reg  [3:0]          reg_pipe5_map6_aggr_id;            
reg  [3:0]          reg_pipe5_map7_aggr_id;            
reg  [3:0]          reg_pipe5_map8_aggr_id;            
reg  [3:0]          reg_pipe5_map9_aggr_id;            
reg  [3:0]          reg_pipe5_map10_aggr_id;            
reg  [3:0]          reg_pipe5_map11_aggr_id;            
reg  [3:0]          reg_pipe5_map12_aggr_id;            
reg  [3:0]          reg_pipe5_map13_aggr_id;            
reg  [3:0]          reg_pipe5_map14_aggr_id;            
reg  [3:0]          reg_pipe5_map15_aggr_id;            
reg  [1:0]          reg_pipe5_map0_vc_source;            
reg  [1:0]          reg_pipe5_map1_vc_source;            
reg  [1:0]          reg_pipe5_map2_vc_source;            
reg  [1:0]          reg_pipe5_map3_vc_source;            
reg  [1:0]          reg_pipe5_map4_vc_source;            
reg  [1:0]          reg_pipe5_map5_vc_source;            
reg  [1:0]          reg_pipe5_map6_vc_source;            
reg  [1:0]          reg_pipe5_map7_vc_source;            
reg  [1:0]          reg_pipe5_map8_vc_source;            
reg  [1:0]          reg_pipe5_map9_vc_source;            
reg  [1:0]          reg_pipe5_map10_vc_source;            
reg  [1:0]          reg_pipe5_map11_vc_source;            
reg  [1:0]          reg_pipe5_map12_vc_source;            
reg  [1:0]          reg_pipe5_map13_vc_source;            
reg  [1:0]          reg_pipe5_map14_vc_source;            
reg  [1:0]          reg_pipe5_map15_vc_source;            
reg  [1:0]          reg_pipe5_map0_vc_dest;            
reg  [1:0]          reg_pipe5_map1_vc_dest;            
reg  [1:0]          reg_pipe5_map2_vc_dest;            
reg  [1:0]          reg_pipe5_map3_vc_dest;            
reg  [1:0]          reg_pipe5_map4_vc_dest;            
reg  [1:0]          reg_pipe5_map5_vc_dest;            
reg  [1:0]          reg_pipe5_map6_vc_dest;            
reg  [1:0]          reg_pipe5_map7_vc_dest;            
reg  [1:0]          reg_pipe5_map8_vc_dest;            
reg  [1:0]          reg_pipe5_map9_vc_dest;            
reg  [1:0]          reg_pipe5_map10_vc_dest;            
reg  [1:0]          reg_pipe5_map11_vc_dest;            
reg  [1:0]          reg_pipe5_map12_vc_dest;            
reg  [1:0]          reg_pipe5_map13_vc_dest;            
reg  [1:0]          reg_pipe5_map14_vc_dest;            
reg  [1:0]          reg_pipe5_map15_vc_dest;            
reg  [5:0]          reg_pipe5_map0_dt_source;            
reg  [5:0]          reg_pipe5_map1_dt_source;            
reg  [5:0]          reg_pipe5_map2_dt_source;            
reg  [5:0]          reg_pipe5_map3_dt_source;            
reg  [5:0]          reg_pipe5_map4_dt_source;            
reg  [5:0]          reg_pipe5_map5_dt_source;            
reg  [5:0]          reg_pipe5_map6_dt_source;            
reg  [5:0]          reg_pipe5_map7_dt_source;            
reg  [5:0]          reg_pipe5_map8_dt_source;            
reg  [5:0]          reg_pipe5_map9_dt_source;            
reg  [5:0]          reg_pipe5_map10_dt_source;            
reg  [5:0]          reg_pipe5_map11_dt_source;            
reg  [5:0]          reg_pipe5_map12_dt_source;            
reg  [5:0]          reg_pipe5_map13_dt_source;            
reg  [5:0]          reg_pipe5_map14_dt_source;            
reg  [5:0]          reg_pipe5_map15_dt_source;            
reg  [5:0]          reg_pipe5_map0_dt_dest;            
reg  [5:0]          reg_pipe5_map1_dt_dest;            
reg  [5:0]          reg_pipe5_map2_dt_dest;            
reg  [5:0]          reg_pipe5_map3_dt_dest;            
reg  [5:0]          reg_pipe5_map4_dt_dest;            
reg  [5:0]          reg_pipe5_map5_dt_dest;            
reg  [5:0]          reg_pipe5_map6_dt_dest;            
reg  [5:0]          reg_pipe5_map7_dt_dest;            
reg  [5:0]          reg_pipe5_map8_dt_dest;            
reg  [5:0]          reg_pipe5_map9_dt_dest;            
reg  [5:0]          reg_pipe5_map10_dt_dest;            
reg  [5:0]          reg_pipe5_map11_dt_dest;            
reg  [5:0]          reg_pipe5_map12_dt_dest;            
reg  [5:0]          reg_pipe5_map13_dt_dest;            
reg  [5:0]          reg_pipe5_map14_dt_dest;            
reg  [5:0]          reg_pipe5_map15_dt_dest;            
reg  [1:0]          reg_pipe5_wr_mode;
wire [31:0]         reg_rd_app_full_cnt_async_fifo_pipe5;
wire [31:0]         reg_rd_app_full_cnt_sync_fifo_pipe5;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_pf_pipe5;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_ph_pipe5;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fe_pipe5;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fs_pipe5;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_le_pipe5;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_ls_pipe5;
reg                reg_clear_app_full_cnt_async_fifo_pipe5;
reg                reg_clear_app_full_cnt_sync_fifo_pipe5;
reg                reg_clear_resv_pkt_cnt_lp_pf_pipe5 ;
reg                reg_clear_resv_pkt_cnt_lp_ph_pipe5 ;
reg                reg_clear_resv_pkt_cnt_sp_fe_pipe5 ;
reg                reg_clear_resv_pkt_cnt_sp_fs_pipe5 ;
reg                reg_clear_resv_pkt_cnt_sp_le_pipe5 ;
reg                reg_clear_resv_pkt_cnt_sp_ls_pipe5 ;
reg                 fifo_wrclk6;
reg                 fifo_rdclk6;
reg                 fifo_wrclk_rst_n6;
reg                 fifo_rdclk_rst_n6;
reg                 reg_line_delay_en6;
reg [1:0]           reg_pipe6_stream_sel;
reg [16:0]          reg_time_window6;
reg                 reg_video_loss_en6;
reg  [15:0]         reg_pipe6_map_en;            
reg  [3:0]          reg_pipe6_map0_aggr_id;            
reg  [3:0]          reg_pipe6_map1_aggr_id;            
reg  [3:0]          reg_pipe6_map2_aggr_id;            
reg  [3:0]          reg_pipe6_map3_aggr_id;            
reg  [3:0]          reg_pipe6_map4_aggr_id;            
reg  [3:0]          reg_pipe6_map5_aggr_id;            
reg  [3:0]          reg_pipe6_map6_aggr_id;            
reg  [3:0]          reg_pipe6_map7_aggr_id;            
reg  [3:0]          reg_pipe6_map8_aggr_id;            
reg  [3:0]          reg_pipe6_map9_aggr_id;            
reg  [3:0]          reg_pipe6_map10_aggr_id;            
reg  [3:0]          reg_pipe6_map11_aggr_id;            
reg  [3:0]          reg_pipe6_map12_aggr_id;            
reg  [3:0]          reg_pipe6_map13_aggr_id;            
reg  [3:0]          reg_pipe6_map14_aggr_id;            
reg  [3:0]          reg_pipe6_map15_aggr_id;            
reg  [1:0]          reg_pipe6_map0_vc_source;            
reg  [1:0]          reg_pipe6_map1_vc_source;            
reg  [1:0]          reg_pipe6_map2_vc_source;            
reg  [1:0]          reg_pipe6_map3_vc_source;            
reg  [1:0]          reg_pipe6_map4_vc_source;            
reg  [1:0]          reg_pipe6_map5_vc_source;            
reg  [1:0]          reg_pipe6_map6_vc_source;            
reg  [1:0]          reg_pipe6_map7_vc_source;            
reg  [1:0]          reg_pipe6_map8_vc_source;            
reg  [1:0]          reg_pipe6_map9_vc_source;            
reg  [1:0]          reg_pipe6_map10_vc_source;            
reg  [1:0]          reg_pipe6_map11_vc_source;            
reg  [1:0]          reg_pipe6_map12_vc_source;            
reg  [1:0]          reg_pipe6_map13_vc_source;            
reg  [1:0]          reg_pipe6_map14_vc_source;            
reg  [1:0]          reg_pipe6_map15_vc_source;            
reg  [1:0]          reg_pipe6_map0_vc_dest;            
reg  [1:0]          reg_pipe6_map1_vc_dest;            
reg  [1:0]          reg_pipe6_map2_vc_dest;            
reg  [1:0]          reg_pipe6_map3_vc_dest;            
reg  [1:0]          reg_pipe6_map4_vc_dest;            
reg  [1:0]          reg_pipe6_map5_vc_dest;            
reg  [1:0]          reg_pipe6_map6_vc_dest;            
reg  [1:0]          reg_pipe6_map7_vc_dest;            
reg  [1:0]          reg_pipe6_map8_vc_dest;            
reg  [1:0]          reg_pipe6_map9_vc_dest;            
reg  [1:0]          reg_pipe6_map10_vc_dest;            
reg  [1:0]          reg_pipe6_map11_vc_dest;            
reg  [1:0]          reg_pipe6_map12_vc_dest;            
reg  [1:0]          reg_pipe6_map13_vc_dest;            
reg  [1:0]          reg_pipe6_map14_vc_dest;            
reg  [1:0]          reg_pipe6_map15_vc_dest;            
reg  [5:0]          reg_pipe6_map0_dt_source;            
reg  [5:0]          reg_pipe6_map1_dt_source;            
reg  [5:0]          reg_pipe6_map2_dt_source;            
reg  [5:0]          reg_pipe6_map3_dt_source;            
reg  [5:0]          reg_pipe6_map4_dt_source;            
reg  [5:0]          reg_pipe6_map5_dt_source;            
reg  [5:0]          reg_pipe6_map6_dt_source;            
reg  [5:0]          reg_pipe6_map7_dt_source;            
reg  [5:0]          reg_pipe6_map8_dt_source;            
reg  [5:0]          reg_pipe6_map9_dt_source;            
reg  [5:0]          reg_pipe6_map10_dt_source;            
reg  [5:0]          reg_pipe6_map11_dt_source;            
reg  [5:0]          reg_pipe6_map12_dt_source;            
reg  [5:0]          reg_pipe6_map13_dt_source;            
reg  [5:0]          reg_pipe6_map14_dt_source;            
reg  [5:0]          reg_pipe6_map15_dt_source;            
reg  [5:0]          reg_pipe6_map0_dt_dest;            
reg  [5:0]          reg_pipe6_map1_dt_dest;            
reg  [5:0]          reg_pipe6_map2_dt_dest;            
reg  [5:0]          reg_pipe6_map3_dt_dest;            
reg  [5:0]          reg_pipe6_map4_dt_dest;            
reg  [5:0]          reg_pipe6_map5_dt_dest;            
reg  [5:0]          reg_pipe6_map6_dt_dest;            
reg  [5:0]          reg_pipe6_map7_dt_dest;            
reg  [5:0]          reg_pipe6_map8_dt_dest;            
reg  [5:0]          reg_pipe6_map9_dt_dest;            
reg  [5:0]          reg_pipe6_map10_dt_dest;            
reg  [5:0]          reg_pipe6_map11_dt_dest;            
reg  [5:0]          reg_pipe6_map12_dt_dest;            
reg  [5:0]          reg_pipe6_map13_dt_dest;            
reg  [5:0]          reg_pipe6_map14_dt_dest;            
reg  [5:0]          reg_pipe6_map15_dt_dest;            
reg  [1:0]          reg_pipe6_wr_mode;
wire [31:0]         reg_rd_app_full_cnt_async_fifo_pipe6;
wire [31:0]         reg_rd_app_full_cnt_sync_fifo_pipe6;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_pf_pipe6;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_ph_pipe6;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fe_pipe6;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fs_pipe6;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_le_pipe6;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_ls_pipe6;
reg                reg_clear_app_full_cnt_async_fifo_pipe6;
reg                reg_clear_app_full_cnt_sync_fifo_pipe6;
reg                reg_clear_resv_pkt_cnt_lp_pf_pipe6 ;
reg                reg_clear_resv_pkt_cnt_lp_ph_pipe6 ;
reg                reg_clear_resv_pkt_cnt_sp_fe_pipe6 ;
reg                reg_clear_resv_pkt_cnt_sp_fs_pipe6 ;
reg                reg_clear_resv_pkt_cnt_sp_le_pipe6 ;
reg                reg_clear_resv_pkt_cnt_sp_ls_pipe6 ;
reg                 fifo_wrclk7;
reg                 fifo_rdclk7;
reg                 fifo_wrclk_rst_n7;
reg                 fifo_rdclk_rst_n7;
reg                 reg_line_delay_en7;
reg [1:0]           reg_pipe7_stream_sel;
reg [16:0]          reg_time_window7;
reg                 reg_video_loss_en7;
reg  [15:0]         reg_pipe7_map_en;            
reg  [3:0]          reg_pipe7_map0_aggr_id;            
reg  [3:0]          reg_pipe7_map1_aggr_id;            
reg  [3:0]          reg_pipe7_map2_aggr_id;            
reg  [3:0]          reg_pipe7_map3_aggr_id;            
reg  [3:0]          reg_pipe7_map4_aggr_id;            
reg  [3:0]          reg_pipe7_map5_aggr_id;            
reg  [3:0]          reg_pipe7_map6_aggr_id;            
reg  [3:0]          reg_pipe7_map7_aggr_id;            
reg  [3:0]          reg_pipe7_map8_aggr_id;            
reg  [3:0]          reg_pipe7_map9_aggr_id;            
reg  [3:0]          reg_pipe7_map10_aggr_id;            
reg  [3:0]          reg_pipe7_map11_aggr_id;            
reg  [3:0]          reg_pipe7_map12_aggr_id;            
reg  [3:0]          reg_pipe7_map13_aggr_id;            
reg  [3:0]          reg_pipe7_map14_aggr_id;            
reg  [3:0]          reg_pipe7_map15_aggr_id;            
reg  [1:0]          reg_pipe7_map0_vc_source;            
reg  [1:0]          reg_pipe7_map1_vc_source;            
reg  [1:0]          reg_pipe7_map2_vc_source;            
reg  [1:0]          reg_pipe7_map3_vc_source;            
reg  [1:0]          reg_pipe7_map4_vc_source;            
reg  [1:0]          reg_pipe7_map5_vc_source;            
reg  [1:0]          reg_pipe7_map6_vc_source;            
reg  [1:0]          reg_pipe7_map7_vc_source;            
reg  [1:0]          reg_pipe7_map8_vc_source;            
reg  [1:0]          reg_pipe7_map9_vc_source;            
reg  [1:0]          reg_pipe7_map10_vc_source;            
reg  [1:0]          reg_pipe7_map11_vc_source;            
reg  [1:0]          reg_pipe7_map12_vc_source;            
reg  [1:0]          reg_pipe7_map13_vc_source;            
reg  [1:0]          reg_pipe7_map14_vc_source;            
reg  [1:0]          reg_pipe7_map15_vc_source;            
reg  [1:0]          reg_pipe7_map0_vc_dest;            
reg  [1:0]          reg_pipe7_map1_vc_dest;            
reg  [1:0]          reg_pipe7_map2_vc_dest;            
reg  [1:0]          reg_pipe7_map3_vc_dest;            
reg  [1:0]          reg_pipe7_map4_vc_dest;            
reg  [1:0]          reg_pipe7_map5_vc_dest;            
reg  [1:0]          reg_pipe7_map6_vc_dest;            
reg  [1:0]          reg_pipe7_map7_vc_dest;            
reg  [1:0]          reg_pipe7_map8_vc_dest;            
reg  [1:0]          reg_pipe7_map9_vc_dest;            
reg  [1:0]          reg_pipe7_map10_vc_dest;            
reg  [1:0]          reg_pipe7_map11_vc_dest;            
reg  [1:0]          reg_pipe7_map12_vc_dest;            
reg  [1:0]          reg_pipe7_map13_vc_dest;            
reg  [1:0]          reg_pipe7_map14_vc_dest;            
reg  [1:0]          reg_pipe7_map15_vc_dest;            
reg  [5:0]          reg_pipe7_map0_dt_source;            
reg  [5:0]          reg_pipe7_map1_dt_source;            
reg  [5:0]          reg_pipe7_map2_dt_source;            
reg  [5:0]          reg_pipe7_map3_dt_source;            
reg  [5:0]          reg_pipe7_map4_dt_source;            
reg  [5:0]          reg_pipe7_map5_dt_source;            
reg  [5:0]          reg_pipe7_map6_dt_source;            
reg  [5:0]          reg_pipe7_map7_dt_source;            
reg  [5:0]          reg_pipe7_map8_dt_source;            
reg  [5:0]          reg_pipe7_map9_dt_source;            
reg  [5:0]          reg_pipe7_map10_dt_source;            
reg  [5:0]          reg_pipe7_map11_dt_source;            
reg  [5:0]          reg_pipe7_map12_dt_source;            
reg  [5:0]          reg_pipe7_map13_dt_source;            
reg  [5:0]          reg_pipe7_map14_dt_source;            
reg  [5:0]          reg_pipe7_map15_dt_source;            
reg  [5:0]          reg_pipe7_map0_dt_dest;            
reg  [5:0]          reg_pipe7_map1_dt_dest;            
reg  [5:0]          reg_pipe7_map2_dt_dest;            
reg  [5:0]          reg_pipe7_map3_dt_dest;            
reg  [5:0]          reg_pipe7_map4_dt_dest;            
reg  [5:0]          reg_pipe7_map5_dt_dest;            
reg  [5:0]          reg_pipe7_map6_dt_dest;            
reg  [5:0]          reg_pipe7_map7_dt_dest;            
reg  [5:0]          reg_pipe7_map8_dt_dest;            
reg  [5:0]          reg_pipe7_map9_dt_dest;            
reg  [5:0]          reg_pipe7_map10_dt_dest;            
reg  [5:0]          reg_pipe7_map11_dt_dest;            
reg  [5:0]          reg_pipe7_map12_dt_dest;            
reg  [5:0]          reg_pipe7_map13_dt_dest;            
reg  [5:0]          reg_pipe7_map14_dt_dest;            
reg  [5:0]          reg_pipe7_map15_dt_dest;            
reg  [1:0]          reg_pipe7_wr_mode;
reg                 reg_pipe0_drop_ls_le_pkt;
reg                 reg_pipe1_drop_ls_le_pkt;
reg                 reg_pipe2_drop_ls_le_pkt;
reg                 reg_pipe3_drop_ls_le_pkt;
reg                 reg_pipe4_drop_ls_le_pkt;
reg                 reg_pipe5_drop_ls_le_pkt;
reg                 reg_pipe6_drop_ls_le_pkt;
reg                 reg_pipe7_drop_ls_le_pkt;
reg  [7:0]          reg_drop_mapping_fault_pkt;
wire [31:0]         reg_rd_app_full_cnt_async_fifo_pipe7;
wire [31:0]         reg_rd_app_full_cnt_sync_fifo_pipe7;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_pf_pipe7;
wire [31:0]         reg_rd_resv_pkt_cnt_lp_ph_pipe7;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fe_pipe7;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_fs_pipe7;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_le_pipe7;
wire [31:0]         reg_rd_resv_pkt_cnt_sp_ls_pipe7;
wire [31:0]         reg_rd_pipe0_dispatched_cnt_ready_for_sch;
wire [31:0]         reg_rd_pipe1_dispatched_cnt_ready_for_sch;
wire [31:0]         reg_rd_pipe2_dispatched_cnt_ready_for_sch;
wire [31:0]         reg_rd_pipe3_dispatched_cnt_ready_for_sch;
wire [31:0]         reg_rd_pipe4_dispatched_cnt_ready_for_sch;
wire [31:0]         reg_rd_pipe5_dispatched_cnt_ready_for_sch;
wire [31:0]         reg_rd_pipe6_dispatched_cnt_ready_for_sch;
wire [31:0]         reg_rd_pipe7_dispatched_cnt_ready_for_sch;
reg                reg_clear_app_full_cnt_async_fifo_pipe7;
reg                reg_clear_app_full_cnt_sync_fifo_pipe7;
reg                reg_clear_resv_pkt_cnt_lp_pf_pipe7 ;
reg                reg_clear_resv_pkt_cnt_lp_ph_pipe7 ;
reg                reg_clear_resv_pkt_cnt_sp_fe_pipe7 ;
reg                reg_clear_resv_pkt_cnt_sp_fs_pipe7 ;
reg                reg_clear_resv_pkt_cnt_sp_le_pipe7 ;
reg                reg_clear_resv_pkt_cnt_sp_ls_pipe7 ;

reg                 reg_resv_pkt_match_lp_dt_en   ;
reg  [5:0]          reg_resv_pkt_match_lp_dt      ;
reg                 reg_clear_resv_pkt_cnt_lp_pf  ;
reg                 reg_clear_resv_pkt_cnt_lp_ph  ;
reg                 reg_clear_resv_pkt_cnt_sp_fe  ;
reg                 reg_clear_resv_pkt_cnt_sp_fs  ;
reg                 reg_clear_resv_pkt_cnt_sp_le  ;
reg                 reg_clear_resv_pkt_cnt_sp_ls  ;
reg                 reg_send_pkt_match_lp_dt_en   ;
reg  [5:0]          reg_send_pkt_match_lp_dt      ;
reg                 reg_clear_send_pkt_cnt_lp_pf  ;
reg                 reg_clear_send_pkt_cnt_lp_ph  ;
reg                 reg_clear_send_pkt_cnt_sp_fe  ;
reg                 reg_clear_send_pkt_cnt_sp_fs  ;
reg                 reg_clear_send_pkt_cnt_sp_le  ;
reg                 reg_clear_send_pkt_cnt_sp_ls  ;
reg                 reg_app_pkt_crc_gen_dis       ;
reg  [3:0]          reg_app_aggr_idi_crc_chk_en   ;
reg  [7:0]          reg_sram_lcrc_err_oen         ;
reg  [7:0]          reg_video_pipe_en             ;

reg             ppi_clk0;        // to u0_dwc_mipicsi2_device_vpg of dwc_mipicsi2_device_vpg.v
reg             ppi_clk1;        // to u1_dwc_mipicsi2_device_vpg of dwc_mipicsi2_device_vpg.v
reg             ppi_clk2;        // to u2_dwc_mipicsi2_device_vpg of dwc_mipicsi2_device_vpg.v
reg             ppi_clk3;        // to u3_dwc_mipicsi2_device_vpg of dwc_mipicsi2_device_vpg.v
reg            ppi_clkrstz0;        // To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            ppi_clkrstz1;        // To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            ppi_clkrstz2;        // To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            ppi_clkrstz3;        // To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_BK_LINES_RS-1:0] vpg_bk_lines_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_BK_LINES_RS-1:0] vpg_bk_lines_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_BK_LINES_RS-1:0] vpg_bk_lines_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_BK_LINES_RS-1:0] vpg_bk_lines_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_DT_RS-1:0] vpg_dt_qst0;    // To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_DT_RS-1:0] vpg_dt_qst1;    // To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_DT_RS-1:0] vpg_dt_qst2;    // To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_DT_RS-1:0] vpg_dt_qst3;    // To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_en0;        // To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_en1;        // To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_en2;        // To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_en3;        // To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_FRAME_NUM_MODE_RS-1:0] vpg_frame_num_mode_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_FRAME_NUM_MODE_RS-1:0] vpg_frame_num_mode_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_FRAME_NUM_MODE_RS-1:0] vpg_frame_num_mode_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_FRAME_NUM_MODE_RS-1:0] vpg_frame_num_mode_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_HBP_TIME_RS-1:0] vpg_hbp_time_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_HBP_TIME_RS-1:0] vpg_hbp_time_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_HBP_TIME_RS-1:0] vpg_hbp_time_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_HBP_TIME_RS-1:0] vpg_hbp_time_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_header_gen_en_lane0;    // To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_header_gen_en1;    // To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_header_gen_en2;    // To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_header_gen_en3;    // To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_HLINE_TIME_RS-1:0] vpg_hline_time_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_HLINE_TIME_RS-1:0] vpg_hline_time_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_HLINE_TIME_RS-1:0] vpg_hline_time_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_HLINE_TIME_RS-1:0] vpg_hline_time_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_HSA_TIME_RS-1:0] vpg_hsa_time_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_HSA_TIME_RS-1:0] vpg_hsa_time_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_HSA_TIME_RS-1:0] vpg_hsa_time_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_HSA_TIME_RS-1:0] vpg_hsa_time_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg           vpg_hsync_packet_en_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg           vpg_hsync_packet_en_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg           vpg_hsync_packet_en_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg           vpg_hsync_packet_en_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_LINE_NUM_MODE_RS-1:0] vpg_line_num_mode_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_LINE_NUM_MODE_RS-1:0] vpg_line_num_mode_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_LINE_NUM_MODE_RS-1:0] vpg_line_num_mode_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_LINE_NUM_MODE_RS-1:0] vpg_line_num_mode_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_MAX_FRAME_NUM_RS-1:0] vpg_max_frame_num_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_MAX_FRAME_NUM_RS-1:0] vpg_max_frame_num_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_MAX_FRAME_NUM_RS-1:0] vpg_max_frame_num_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_MAX_FRAME_NUM_RS-1:0] vpg_max_frame_num_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_mode_qst0;        // To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_mode_qst1;        // To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_mode_qst2;        // To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_mode_qst3;        // To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_orientation_qst0;    // To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_orientation_qst1;    // To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_orientation_qst2;    // To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_orientation_qst3;    // To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_packet_lost_ack0;    // To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_packet_lost_ack1;    // To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_packet_lost_ack2;    // To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_packet_lost_ack3;    // To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_payload_gen_en0;    // To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_payload_gen_en1;    // To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_payload_gen_en2;    // To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg            vpg_payload_gen_en3;    // To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_PKT_SIZE_RS-1:0] vpg_pkt_size_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_PKT_SIZE_RS-1:0] vpg_pkt_size_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_PKT_SIZE_RS-1:0] vpg_pkt_size_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_PKT_SIZE_RS-1:0] vpg_pkt_size_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_START_LINE_NUM_RS-1:0] vpg_start_line_num_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_START_LINE_NUM_RS-1:0] vpg_start_line_num_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_START_LINE_NUM_RS-1:0] vpg_start_line_num_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_START_LINE_NUM_RS-1:0] vpg_start_line_num_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_STEP_LINE_NUM_RS-1:0] vpg_step_line_num_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_STEP_LINE_NUM_RS-1:0] vpg_step_line_num_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_STEP_LINE_NUM_RS-1:0] vpg_step_line_num_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_STEP_LINE_NUM_RS-1:0] vpg_step_line_num_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_ACT_LINES_RS-1:0] vpg_vactive_lines_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_ACT_LINES_RS-1:0] vpg_vactive_lines_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_ACT_LINES_RS-1:0] vpg_vactive_lines_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_ACT_LINES_RS-1:0] vpg_vactive_lines_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VBP_LINES_RS-1:0] vpg_vbp_lines_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VBP_LINES_RS-1:0] vpg_vbp_lines_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VBP_LINES_RS-1:0] vpg_vbp_lines_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VBP_LINES_RS-1:0] vpg_vbp_lines_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VC_RS-1:0] vpg_vc_qst0;    // To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VC_RS-1:0] vpg_vc_qst1;    // To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VC_RS-1:0] vpg_vc_qst2;    // To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VC_RS-1:0] vpg_vc_qst3;    // To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VCX_DWIDTH-1:0] vpg_vcx_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VCX_DWIDTH-1:0] vpg_vcx_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VCX_DWIDTH-1:0] vpg_vcx_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VCX_DWIDTH-1:0] vpg_vcx_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VFP_LINES_RS-1:0] vpg_vfp_lines_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VFP_LINES_RS-1:0] vpg_vfp_lines_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VFP_LINES_RS-1:0] vpg_vfp_lines_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VFP_LINES_RS-1:0] vpg_vfp_lines_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VSA_LINES_RS-1:0] vpg_vsa_lines_qst0;// To u0_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VSA_LINES_RS-1:0] vpg_vsa_lines_qst1;// To u1_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VSA_LINES_RS-1:0] vpg_vsa_lines_qst2;// To u2_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg [CSI2_DEVICE_VPG_VSA_LINES_RS-1:0] vpg_vsa_lines_qst3;// To u3_DWC_mipicsi2_device_vpg of DWC_mipicsi2_device_vpg.v
reg                                    reg_mipi_host_sel;
/***as6s_app_vprbs_gen,as6s_app_vprbs_chk***/
reg  [15:0]         reg_vprbs_tx_idi_driver_pkt_interval            ;
reg  [15:0]         reg_vprbs_tx_idi_driver_total_interval          ;
reg  [5:0]          reg_vprbs_tx_idi_driver_data_type               ;
reg  [3:0]          reg_vprbs_tx_idi_driver_virtual_channel         ;
reg  [15:0]         reg_vprbs_tx_idi_driver_word_count              ;
reg                 reg_vprbs_tx_err_inject_en                      ;
reg  [7:0]          reg_vprbs_tx_err_inject_intv_num                ;
reg  [7:0]          reg_vprbs_tx_err_inject_intv_time               ;
reg                 reg_vprbs_tx_gen_en                             ;
reg  [2:0]          reg_vprbs_tx_mode                               ;
reg                 reg_vprbs_tx_order                              ;
reg                 reg_vprbs_tx_pat_reset                          ;
reg                 reg_vprbs_loopback                              ;
reg                 reg_vprbs_rx_chk_en                             ;
reg  [2:0]          reg_vprbs_rx_mode                               ;
reg                 reg_vprbs_rx_order                              ;
reg                 reg_vprbs_rx_load                               ;
reg                 reg_vprbs_rx_lock_continue                      ;
reg  [3:0]          reg_vprbs_rx_locked_match_cnt                   ;
reg  [3:0]          reg_vprbs_rx_uncheck_tolerance                  ;
reg                 reg_vprbs_rx_err_clear                          ;
reg                 reg_sch0_fse_filter                             ;
reg                 reg_sch1_fse_filter                             ;
reg                 reg_sch2_fse_filter                             ;
reg                 reg_sch3_fse_filter                             ;
reg                 reg_app_wr_idi_data_continue                    ;


wire                dvp_afifo_ovf_int;
wire                dvp_afifo_udf_int;
wire    [15:0]      idi_vpg_word_count_lane0;
wire    [2 :0]      idi_vpg_byte_en_lane0;
wire                idi_vpg_header_en_lane0;
wire                idi_vpg_data_en_lane0;
wire    [63:0]      idi_vpg_data_lane0;
wire    [1 :0]      idi_vpg_vc_lane0;
wire    [1 :0]      idi_vpg_vcx_lane0;
wire    [5 :0]      idi_vpg_dt_lane0;
wire    [15:0]      idi_vpg_word_count_lane1;
wire    [2 :0]      idi_vpg_byte_en_lane1;
wire                idi_vpg_header_en_lane1;
wire                idi_vpg_data_en_lane1;
wire    [63:0]      idi_vpg_data_lane1;
wire    [1 :0]      idi_vpg_vc_lane1;
wire    [1 :0]      idi_vpg_vcx_lane1;
wire    [5 :0]      idi_vpg_dt_lane1;
wire    [15:0]      idi_vpg_word_count_lane2;
wire    [2 :0]      idi_vpg_byte_en_lane2;
wire                idi_vpg_header_en_lane2;
wire                idi_vpg_data_en_lane2;
wire    [63:0]      idi_vpg_data_lane2;
wire    [1 :0]      idi_vpg_vc_lane2;
wire    [1 :0]      idi_vpg_vcx_lane2;
wire    [5 :0]      idi_vpg_dt_lane2;
wire    [15:0]      idi_vpg_word_count_lane3;
wire    [2 :0]      idi_vpg_byte_en_lane3;
wire                idi_vpg_header_en_lane3;
wire                idi_vpg_data_en_lane3;
wire    [63:0]      idi_vpg_data_lane3;
wire    [1 :0]      idi_vpg_vc_lane3;
wire    [1 :0]      idi_vpg_vcx_lane3;
wire    [5 :0]      idi_vpg_dt_lane3;

wire    [15:0]      idi_word_count_lane0;
wire    [2 :0]      idi_byte_en_lane0;
wire                idi_header_en_lane0;
wire                idi_data_en_lane0;
wire    [63:0]      idi_data_lane0;
wire    [1 :0]      idi_vc_lane0;
wire    [1 :0]      idi_vcx_lane0;
wire    [5 :0]      idi_dt_lane0;
wire    [15:0]      idi_word_count_lane1;
wire    [2 :0]      idi_byte_en_lane1;
wire                idi_header_en_lane1;
wire                idi_data_en_lane1;
wire    [63:0]      idi_data_lane1;
wire    [1 :0]      idi_vc_lane1;
wire    [1 :0]      idi_vcx_lane1;
wire    [5 :0]      idi_dt_lane1;
wire    [15:0]      idi_word_count_lane2;
wire    [2 :0]      idi_byte_en_lane2;
wire                idi_header_en_lane2;
wire                idi_data_en_lane2;
wire    [63:0]      idi_data_lane2;
wire    [1 :0]      idi_vc_lane2;
wire    [1 :0]      idi_vcx_lane2;
wire    [5 :0]      idi_dt_lane2;
wire    [15:0]      idi_word_count_lane3;
wire    [2 :0]      idi_byte_en_lane3;
wire                idi_header_en_lane3;
wire                idi_data_en_lane3;
wire    [63:0]      idi_data_lane3;
wire    [1 :0]      idi_vc_lane3;
wire    [1 :0]      idi_vcx_lane3;
wire    [5 :0]      idi_dt_lane3;

reg                 app_clk_data;        
reg                 app_clk_rst_n;        

wire    [3:0]       idi_prbs_chk_byte_en            ;
wire    [127:0]     idi_prbs_chk_data               ;
wire                idi_prbs_chk_data_en            ;
wire    [20:0]      idi_prbs_chk_data_parity        ;
wire    [5:0]       idi_prbs_chk_data_type          ;
wire                idi_prbs_chk_header_en          ;
wire    [1:0]       idi_prbs_chk_virtual_channel    ;
wire    [2:0]       idi_prbs_chk_virtual_channel_x  ;
wire    [15:0]      idi_prbs_chk_word_count         ;

reg			    reg_vprbs_rx_chk_en0            ;
reg			    reg_vprbs_rx_chk_en1            ;
reg			    reg_vprbs_rx_chk_en2            ;
reg			    reg_vprbs_rx_chk_en3            ;
reg			    reg_vprbs_rx_chk_en4            ;
reg			    reg_vprbs_rx_chk_en5            ;
reg			    reg_vprbs_rx_chk_en6            ;
reg			    reg_vprbs_rx_chk_en7            ;
reg			    reg_vprbs_tx_gen_en0            ;
reg			    reg_vprbs_tx_gen_en1            ;
reg			    reg_vprbs_tx_gen_en2            ;
reg			    reg_vprbs_tx_gen_en3            ;
reg			    reg_vprbs_tx_gen_en4            ;
reg			    reg_vprbs_tx_gen_en5            ;
reg			    reg_vprbs_tx_gen_en6            ;
reg			    reg_vprbs_tx_gen_en7            ;
wire            reg_dvp_mode_en                 ;
reg             reg_dvp_mode_en_bank2app        ;
reg			    reg_dbl_mode;
reg [4:0]		reg_crossbar_0;
reg [4:0]		reg_crossbar_1;
reg [4:0]		reg_crossbar_10;
reg [4:0]		reg_crossbar_11;
reg [4:0]		reg_crossbar_12;
reg [4:0]		reg_crossbar_13;
reg [4:0]		reg_crossbar_14;
reg [4:0]		reg_crossbar_15;
reg [4:0]		reg_crossbar_16;
reg [4:0]		reg_crossbar_17;
reg [4:0]		reg_crossbar_18;
reg [4:0]		reg_crossbar_19;
reg [4:0]		reg_crossbar_2;
reg [4:0]		reg_crossbar_20;
reg [4:0]		reg_crossbar_21;
reg [4:0]		reg_crossbar_22;
reg [4:0]		reg_crossbar_23;
reg [4:0]		reg_crossbar_3;
reg [4:0]		reg_crossbar_4;
reg [4:0]		reg_crossbar_5;
reg [4:0]		reg_crossbar_6;
reg [4:0]		reg_crossbar_7;
reg [4:0]		reg_crossbar_8;
reg [4:0]		reg_crossbar_9;
reg [4:0]		reg_crossbar_vs;
reg [4:0]		reg_crossbar_hs;
reg [31:0]		reg_de_cnt;
reg [31:0]		reg_de_high;
reg [31:0]		reg_de_low;
reg	[5:0]       reg_force_dvp_data_type;
reg	[3:0]	    reg_force_dvp_virtual_channel;
reg	[15:0]	    reg_force_dvp_word_count;
reg             reg_force_dvp_word_count_en;
reg			    reg_force_mux_0;
reg			    reg_force_mux_1;
reg			    reg_force_mux_10;
reg			    reg_force_mux_11;
reg			    reg_force_mux_12;
reg			    reg_force_mux_13;
reg			    reg_force_mux_14;
reg			    reg_force_mux_15;
reg			    reg_force_mux_16;
reg			    reg_force_mux_17;
reg			    reg_force_mux_18;
reg			    reg_force_mux_19;
reg			    reg_force_mux_2;
reg			    reg_force_mux_20;
reg			    reg_force_mux_21;
reg			    reg_force_mux_22;
reg			    reg_force_mux_23;
reg			    reg_force_mux_3;
reg			    reg_force_mux_4;
reg			    reg_force_mux_5;
reg			    reg_force_mux_6;
reg			    reg_force_mux_7;
reg			    reg_force_mux_8;
reg			    reg_force_mux_9;
reg			    reg_force_mux_vs;
reg			    reg_force_mux_hs;
reg			    reg_invert_mux_0;
reg			    reg_invert_mux_1;
reg			    reg_invert_mux_10;
reg			    reg_invert_mux_11;
reg			    reg_invert_mux_12;
reg			    reg_invert_mux_13;
reg			    reg_invert_mux_14;
reg			    reg_invert_mux_15;
reg			    reg_invert_mux_16;
reg			    reg_invert_mux_17;
reg			    reg_invert_mux_18;
reg			    reg_invert_mux_19;
reg			    reg_invert_mux_2;
reg			    reg_invert_mux_20;
reg			    reg_invert_mux_21;
reg			    reg_invert_mux_22;
reg			    reg_invert_mux_23;
reg			    reg_invert_mux_3;
reg			    reg_invert_mux_4;
reg			    reg_invert_mux_5;
reg			    reg_invert_mux_6;
reg			    reg_invert_mux_7;
reg			    reg_invert_mux_8;
reg			    reg_invert_mux_9;
reg			    reg_invert_mux_vs;
reg			    reg_invert_mux_hs;
reg [31:0]		reg_vs2de_dly;
reg [31:0]		reg_vs2fe_dly;
reg [31:0]		reg_vs2fs_dly;
reg [31:0]		reg_hs2de_dly;
reg             reg_vs2de_trigger_en;
reg             reg_hs2de_trigger_en;
reg             reg_dvp_test_en;
reg [15:0]      reg_frame_delay;
reg [15:0]      reg_total_h;
reg [15:0]      reg_total_v;
reg [15:0]      reg_col_start;
reg [15:0]      reg_col_end;
reg [15:0]      reg_row_start;
reg [15:0]      reg_row_end;
reg [15:0]      reg_col_start_hsync_pre_high;
reg [5:0]       reg_data_type;
wire[13:0]      pixel_data;
wire            vsync;
reg             reg_yuyv_mode_en;
wire [15:0]     reg_rd_dvp_clk_cnt_at_clk_10K;
wire [15:0]     reg_rd_dvp_pin_square_det_succeed;
reg             reg_dvp_clk_frequence_det_en;
reg             reg_dvp_pin_square_det_en;
reg             reg_dvp_trigger_en;
reg             reg_dvp_vprbs_tx_gen_en;
reg  [2:0]      reg_dvp_vprbs_tx_mode;
reg             reg_dvp_vprbs_tx_order;
reg  [15:0]     reg_dvp_vprbs_tx_vs_interval;
reg             efuse_filedname_valid;
reg             efuse_info_mipi_en;

wire [2:0]      as6s_csi_bytes_en;
wire [63:0]     as6s_csi_data;
wire			as6s_csi_data_en;
wire [5:0]		as6s_csi_data_type;
wire			as6s_csi_header_en;
reg             reg_video_data_fwft_fifo_ovf_int_mask0;
reg             reg_video_data_fwft_fifo_ovf_int_mask1;
reg             reg_video_data_fwft_fifo_ovf_int_mask2;
reg             reg_video_data_fwft_fifo_ovf_int_mask3;
reg             reg_video_data_fwft_fifo_ovf_int_mask4;
reg             reg_video_data_fwft_fifo_ovf_int_mask5;
reg             reg_video_data_fwft_fifo_ovf_int_mask6;
reg             reg_video_data_fwft_fifo_ovf_int_mask7;
reg             reg_sch0_frame_sync_auto_change_pipe_wr_mode;
reg             reg_sch1_frame_sync_auto_change_pipe_wr_mode;
reg             reg_sch2_frame_sync_auto_change_pipe_wr_mode;
reg             reg_sch3_frame_sync_auto_change_pipe_wr_mode;

initial begin
    efuse_filedname_valid   = 1'd0;
    efuse_info_mipi_en      = 1'd0;
    clk_1M_rst_n        = 1'd0;
    dvp_clk_rst_n       = 1'd0;
    ppi_clkrstz0        = 1'd0;        
    ppi_clkrstz1        = 1'd0;        
    ppi_clkrstz2        = 1'd0;        
    ppi_clkrstz3        = 1'd0;        
    aggre_clk_rst_n0    = 1'd0;    
    aggre_clk_rst_n1    = 1'd0;    
    aggre_clk_rst_n2    = 1'd0;    
    aggre_clk_rst_n3    = 1'd0;    
    fifo_wrclk_rst_n0   = 1'd0;    
    fifo_wrclk_rst_n1   = 1'd0;    
    fifo_wrclk_rst_n2   = 1'd0;    
    fifo_wrclk_rst_n3   = 1'd0;    
    fifo_wrclk_rst_n4   = 1'd0;    
    fifo_wrclk_rst_n5   = 1'd0;    
    fifo_wrclk_rst_n6   = 1'd0;    
    fifo_wrclk_rst_n7   = 1'd0;    
    fifo_rdclk_rst_n0   = 1'd0;    
    fifo_rdclk_rst_n1   = 1'd0;    
    fifo_rdclk_rst_n2   = 1'd0;    
    fifo_rdclk_rst_n3   = 1'd0;    
    fifo_rdclk_rst_n4   = 1'd0;    
    fifo_rdclk_rst_n5   = 1'd0;    
    fifo_rdclk_rst_n6   = 1'd0;    
    fifo_rdclk_rst_n7   = 1'd0;    
    app_clk_rst_n       = 1'd0;
    treed_reg_bank_clk_reset_n  =   1'd0;
    vpg_en0             = 1'd0;
    vpg_en1             = 1'd0;
    vpg_en2             = 1'd0;
    vpg_en3             = 1'd0;
    reg_pipe_fifo_full_clear                    =   4'd0;
    reg_pipe_fifo_full_clear_last_four          =   4'd0;


    #100    
    clk_1M_rst_n        = 1'd1;
    dvp_clk_rst_n       = 1'd1;
    ppi_clkrstz0        = 1'd1;        
    ppi_clkrstz1        = 1'd1;        
    ppi_clkrstz2        = 1'd1;        
    ppi_clkrstz3        = 1'd1;        
    aggre_clk_rst_n0    = 1'd1;    
    aggre_clk_rst_n1    = 1'd1;    
    aggre_clk_rst_n2    = 1'd1;    
    aggre_clk_rst_n3    = 1'd1;    
    fifo_wrclk_rst_n0   = 1'd1;    
    fifo_wrclk_rst_n1   = 1'd1;    
    fifo_wrclk_rst_n2   = 1'd1;    
    fifo_wrclk_rst_n3   = 1'd1;    
    fifo_wrclk_rst_n4   = 1'd1;    
    fifo_wrclk_rst_n5   = 1'd1;    
    fifo_wrclk_rst_n6   = 1'd1;    
    fifo_wrclk_rst_n7   = 1'd1;    
    fifo_rdclk_rst_n0   = 1'd1;    
    fifo_rdclk_rst_n1   = 1'd1;    
    fifo_rdclk_rst_n2   = 1'd1;    
    fifo_rdclk_rst_n3   = 1'd1;    
    fifo_rdclk_rst_n4   = 1'd1;    
    fifo_rdclk_rst_n5   = 1'd1;    
    fifo_rdclk_rst_n6   = 1'd1;    
    fifo_rdclk_rst_n7   = 1'd1;    
    app_clk_rst_n       = 1'd1;
    treed_reg_bank_clk_reset_n  =   1'd1;
    #100
    vpg_en0             = 1'd1;
    vpg_en1             = 1'd1;
    vpg_en2             = 1'd1;
    vpg_en3             = 1'd1;

    @(posedge fifo_wrclk0);
    @(posedge fifo_wrclk1);
    @(posedge fifo_wrclk2);
    @(posedge fifo_wrclk3);
    @(posedge fifo_wrclk4);
    @(posedge fifo_wrclk5);
    @(posedge fifo_wrclk6);
    @(posedge fifo_wrclk7);
    reg_pipe0_wr_mode           =   2'b11           ;
    reg_pipe1_wr_mode           =   2'b11           ;
    reg_pipe2_wr_mode           =   2'b11           ;
    reg_pipe3_wr_mode           =   2'b11           ;
    reg_pipe4_wr_mode           =   2'b11           ;
    reg_pipe5_wr_mode           =   2'b11           ;
    reg_pipe6_wr_mode           =   2'b11           ;
    reg_pipe7_wr_mode           =   2'b11           ;
    reg_all_pipe_wr_mode_strobe =   1'd1            ;
    @(posedge fifo_wrclk0);
    @(posedge fifo_wrclk1);
    @(posedge fifo_wrclk2);
    @(posedge fifo_wrclk3);
    @(posedge fifo_wrclk4);
    @(posedge fifo_wrclk5);
    @(posedge fifo_wrclk6);
    @(posedge fifo_wrclk7);
    reg_all_pipe_wr_mode_strobe =   1'd0            ;

    #100
    dvp_clk_rst_n       = 1'd1;
    reg_vprbs_rx_chk_en0  = 1'd1 ;
    reg_vprbs_rx_chk_en1  = 1'd1 ;
    reg_vprbs_rx_chk_en2  = 1'd1 ;
    reg_vprbs_rx_chk_en3  = 1'd1 ;
    reg_vprbs_rx_chk_en4  = 1'd1 ;
    reg_vprbs_rx_chk_en5  = 1'd1 ;
    reg_vprbs_rx_chk_en6  = 1'd1 ;
    reg_vprbs_rx_chk_en7  = 1'd1 ;
    reg_vprbs_tx_gen_en0  = 1'd1 ;
    reg_vprbs_tx_gen_en1  = 1'd1 ;
    reg_vprbs_tx_gen_en2  = 1'd1 ;
    reg_vprbs_tx_gen_en3  = 1'd1 ;
    reg_vprbs_tx_gen_en4  = 1'd1 ;
    reg_vprbs_tx_gen_en5  = 1'd1 ;
    reg_vprbs_tx_gen_en6  = 1'd1 ;
    reg_vprbs_tx_gen_en7  = 1'd1 ;

    #200
	reg_dvp_test_en                 = 1'd1;        

    #1ms
    vpg_en0             = 1'd0;
    vpg_en1             = 1'd0;
    vpg_en2             = 1'd0;
    vpg_en3             = 1'd1;
end



wire[7:0]    idi_ecc_lane0            ;
wire[15:0]    idi_dvalid_lane0        ;
wire[15:0]    idi_hvalid_lane0        ;
wire[15:0]    idi_vvalid_lane0        ;
assign    idi_ecc_lane0                =8'd0;    
assign    idi_dvalid_lane0            =`MEP_CSI2_HOST_N_VIRT_CH'd0;
assign    idi_hvalid_lane0            =`MEP_CSI2_HOST_N_VIRT_CH'd0;
assign    idi_vvalid_lane0            =`MEP_CSI2_HOST_N_VIRT_CH'd0;

initial begin
    reg_video_data_fwft_fifo_ovf_int_mask0  =   1'd0;
    reg_video_data_fwft_fifo_ovf_int_mask1  =   1'd0;
    reg_video_data_fwft_fifo_ovf_int_mask2  =   1'd0;
    reg_video_data_fwft_fifo_ovf_int_mask3  =   1'd0;
    reg_video_data_fwft_fifo_ovf_int_mask4  =   1'd0;
    reg_video_data_fwft_fifo_ovf_int_mask5  =   1'd0;
    reg_video_data_fwft_fifo_ovf_int_mask6  =   1'd0;
    reg_video_data_fwft_fifo_ovf_int_mask7  =   1'd0;
	//reg_vprbs_tx_idi_driver_pkt_interval    =   16'd20          ;
	//reg_vprbs_tx_idi_driver_total_interval  =   16'd100         ;
	//reg_vprbs_tx_idi_driver_data_type       =   6'h24           ;
	//reg_vprbs_tx_idi_driver_virtual_channel =   4'd0            ;
	//reg_vprbs_tx_idi_driver_word_count      =   16'd708         ;
	reg_vprbs_tx_idi_driver_pkt_interval    =   16'd10          ;
	reg_vprbs_tx_idi_driver_total_interval  =   16'd200         ;
	reg_vprbs_tx_idi_driver_data_type       =   6'h24           ;
	reg_vprbs_tx_idi_driver_virtual_channel =   4'd0            ;
	reg_vprbs_tx_idi_driver_word_count      =   16'd3072         ;
    reg_vprbs_tx_err_inject_en              =   1'd1            ;
    reg_vprbs_tx_err_inject_intv_num        =   8'd1            ;
    reg_vprbs_tx_err_inject_intv_time       =   8'd10           ;
    reg_vprbs_tx_gen_en                     =   1'd0            ;
    reg_vprbs_tx_mode                       =   3'd0            ;
    reg_vprbs_tx_order                      =   1'd0            ;
    reg_vprbs_tx_pat_reset                  =   1'd0            ;
    reg_vprbs_loopback                      =   1'd0            ;
    reg_vprbs_rx_chk_en                     =   1'd1            ;
    reg_vprbs_rx_mode                       =   3'd0            ;
    reg_vprbs_rx_order                      =   1'd0            ;
    reg_vprbs_rx_load                       =   1'd1            ;
    reg_vprbs_rx_lock_continue              =   1'd1            ;
    reg_vprbs_rx_locked_match_cnt           =   4'd1            ;
    reg_vprbs_rx_uncheck_tolerance          =   4'd1            ;
    reg_vprbs_rx_err_clear                  =   1'd0            ;
    reg_dvp_trigger_en                      =   1'd1            ;
    reg_dvp_clk_frequence_det_en            =   1'd0            ;
    reg_dvp_pin_square_det_en               =   1'd0            ;
    reg_dvp_vprbs_tx_gen_en                 =   1'd0            ;
    reg_dvp_vprbs_tx_mode                   =   3'd0            ;
    reg_dvp_vprbs_tx_order                  =   1'd0            ;
    reg_dvp_vprbs_tx_vs_interval            =   16'd1000        ; 
    reg_hs2de_dly                           =   32'd1000        ;
    reg_vs2de_trigger_en                    =   1'd1            ;
    reg_dvp_trigger_en                      =   1'd1            ;
    reg_col_start_hsync_pre_high            =   1'd1            ;
end

/*  dvp_driver  AUTO_TEMPLATE (
    .clk(app_clk_data),
    .rst_n(app_clk_rst_n),
)*/
dvp_driver u_dvp_driver(/*AUTOINST*/
			// Outputs
			.pixel_vld	(pixel_vld),
			.pixel_data	(pixel_data[13:0]),
			.vsync		(vsync),
			.hsync		(hsync),
			// Inputs
			.clk		(app_clk_data),		 // Templated
			.rst_n		(app_clk_rst_n),	 // Templated
			.reg_dvp_test_en(reg_dvp_test_en),
			.reg_yuyv_mode_en(reg_yuyv_mode_en),
			.reg_frame_delay(reg_frame_delay[15:0]),
			.reg_total_h	(reg_total_h[15:0]),
			.reg_total_v	(reg_total_v[15:0]),
			.reg_col_start	(reg_col_start[15:0]),
			.reg_col_end	(reg_col_end[15:0]),
			.reg_row_start	(reg_row_start[15:0]),
			.reg_row_end	(reg_row_end[15:0]),
			.reg_data_type	(reg_data_type[5:0]),
			.reg_col_start_hsync_pre_high(reg_col_start_hsync_pre_high[15:0]));



/*  pattern_test  AUTO_TEMPLATE (
	.chk_clk		(ppi_clk0),
	.chk_rst_n		(ppi_clkrstz0),
	.gen_clk		(ppi_clk0),
	.gen_rst_n		(ppi_clkrstz0),
    .idi_gen_data_type	(),
    .idi_gen_header_en	(),
    .idi_gen_virtual_channel(),
    .idi_gen_word_count	(),
    .reg_rd_vprbs_rx_check	(),
    .reg_rd_vprbs_rx_err	(),
    .reg_rd_vprbs_rx_fail	(),
    .idi_gen_data	(),
    .idi_gen_byte_en	(),
    .idi_gen_data_en	(),

	.idi_chk_byte_en	(3'd0),
	.idi_chk_data	(64'd0),
	.idi_chk_data_en	(1'd0),
    .idi_chk_header_en	(1'd0),
    .idi_chk_data_type	(6'd0),
)*/
pattern_test u_pattern_test(/*AUTOINST*/
			    // Outputs
			    .idi_gen_virtual_channel(),		 // Templated
			    .idi_gen_word_count	(),		 // Templated
			    .reg_rd_vprbs_rx_check(),		 // Templated
			    .reg_rd_vprbs_rx_err(),		 // Templated
			    .reg_rd_vprbs_rx_fail(),		 // Templated
			    .idi_gen_header_en	(),		 // Templated
			    .idi_gen_data_en	(),		 // Templated
			    .idi_gen_byte_en	(),		 // Templated
			    .idi_gen_data	(),		 // Templated
			    .idi_gen_data_type	(),		 // Templated
			    // Inputs
			    .chk_clk		(ppi_clk0),	 // Templated
			    .chk_rst_n		(ppi_clkrstz0),	 // Templated
			    .gen_clk		(ppi_clk0),	 // Templated
			    .gen_rst_n		(ppi_clkrstz0),	 // Templated
			    .reg_vprbs_rx_chk_en(reg_vprbs_rx_chk_en),
			    .reg_vprbs_rx_err_clear(reg_vprbs_rx_err_clear),
			    .reg_vprbs_rx_load	(reg_vprbs_rx_load),
			    .reg_vprbs_rx_lock_continue(reg_vprbs_rx_lock_continue),
			    .reg_vprbs_rx_locked_match_cnt(reg_vprbs_rx_locked_match_cnt[3:0]),
			    .reg_vprbs_rx_mode	(reg_vprbs_rx_mode[2:0]),
			    .reg_vprbs_rx_order	(reg_vprbs_rx_order),
			    .reg_vprbs_rx_uncheck_tolerance(reg_vprbs_rx_uncheck_tolerance[3:0]),
			    .reg_vprbs_tx_err_inject_en(reg_vprbs_tx_err_inject_en),
			    .reg_vprbs_tx_err_inject_intv_num(reg_vprbs_tx_err_inject_intv_num[7:0]),
			    .reg_vprbs_tx_err_inject_intv_time(reg_vprbs_tx_err_inject_intv_time[7:0]),
			    .reg_vprbs_tx_gen_en(reg_vprbs_tx_gen_en),
			    .reg_vprbs_tx_idi_driver_data_type(reg_vprbs_tx_idi_driver_data_type[5:0]),
			    .reg_vprbs_tx_idi_driver_pkt_interval(reg_vprbs_tx_idi_driver_pkt_interval[15:0]),
			    .reg_vprbs_tx_idi_driver_total_interval(reg_vprbs_tx_idi_driver_total_interval[15:0]),
			    .reg_vprbs_tx_idi_driver_virtual_channel(reg_vprbs_tx_idi_driver_virtual_channel[3:0]),
			    .reg_vprbs_tx_idi_driver_word_count(reg_vprbs_tx_idi_driver_word_count[15:0]),
			    .reg_vprbs_tx_mode	(reg_vprbs_tx_mode[2:0]),
			    .reg_vprbs_tx_order	(reg_vprbs_tx_order),
			    .reg_vprbs_tx_pat_reset(reg_vprbs_tx_pat_reset),
			    .idi_chk_header_en	(1'd0),		 // Templated
			    .idi_chk_data_en	(1'd0),		 // Templated
			    .idi_chk_byte_en	(3'd0),		 // Templated
			    .idi_chk_data_type	(6'd0),		 // Templated
			    .idi_chk_data	(64'd0),	 // Templated
			    .reg_vprbs_loopback	(reg_vprbs_loopback));

/*  pattern_test  AUTO_TEMPLATE (
	.chk_clk		(app_clk_data),
	.chk_rst_n		(app_clk_rst_n),
	.gen_clk		(app_clk_data),
	.gen_rst_n		(app_clk_rst_n),
    .idi_gen_data_type	(),
    .idi_gen_header_en	(),
    .idi_gen_virtual_channel(),
    .idi_gen_word_count	(),
    .reg_rd_vprbs_rx_check	(),
    .reg_rd_vprbs_rx_err	(),
    .reg_rd_vprbs_rx_fail	(),
    .idi_gen_data	(),
    .idi_gen_byte_en	(),
    .idi_gen_data_en	(),

	.idi_chk_byte_en	(as6s_csi_bytes_en[]),
	.idi_chk_data	    (as6s_csi_data[]),
	.idi_chk_data_en	(as6s_csi_data_en),
    .idi_chk_header_en	(as6s_csi_header_en),
    .idi_chk_data_type	(as6s_csi_data_type[]),
)*/
pattern_test pattern_test_as6s_app_ate(/*AUTOINST*/
				       // Outputs
				       .idi_gen_virtual_channel(),	 // Templated
				       .idi_gen_word_count(),		 // Templated
				       .reg_rd_vprbs_rx_check(),	 // Templated
				       .reg_rd_vprbs_rx_err(),		 // Templated
				       .reg_rd_vprbs_rx_fail(),		 // Templated
				       .idi_gen_header_en(),		 // Templated
				       .idi_gen_data_en	(),		 // Templated
				       .idi_gen_byte_en	(),		 // Templated
				       .idi_gen_data	(),		 // Templated
				       .idi_gen_data_type(),		 // Templated
				       // Inputs
				       .chk_clk		(app_clk_data),	 // Templated
				       .chk_rst_n	(app_clk_rst_n), // Templated
				       .gen_clk		(app_clk_data),	 // Templated
				       .gen_rst_n	(app_clk_rst_n), // Templated
				       .reg_vprbs_rx_chk_en(reg_vprbs_rx_chk_en),
				       .reg_vprbs_rx_err_clear(reg_vprbs_rx_err_clear),
				       .reg_vprbs_rx_load(reg_vprbs_rx_load),
				       .reg_vprbs_rx_lock_continue(reg_vprbs_rx_lock_continue),
				       .reg_vprbs_rx_locked_match_cnt(reg_vprbs_rx_locked_match_cnt[3:0]),
				       .reg_vprbs_rx_mode(reg_vprbs_rx_mode[2:0]),
				       .reg_vprbs_rx_order(reg_vprbs_rx_order),
				       .reg_vprbs_rx_uncheck_tolerance(reg_vprbs_rx_uncheck_tolerance[3:0]),
				       .reg_vprbs_tx_err_inject_en(reg_vprbs_tx_err_inject_en),
				       .reg_vprbs_tx_err_inject_intv_num(reg_vprbs_tx_err_inject_intv_num[7:0]),
				       .reg_vprbs_tx_err_inject_intv_time(reg_vprbs_tx_err_inject_intv_time[7:0]),
				       .reg_vprbs_tx_gen_en(reg_vprbs_tx_gen_en),
				       .reg_vprbs_tx_idi_driver_data_type(reg_vprbs_tx_idi_driver_data_type[5:0]),
				       .reg_vprbs_tx_idi_driver_pkt_interval(reg_vprbs_tx_idi_driver_pkt_interval[15:0]),
				       .reg_vprbs_tx_idi_driver_total_interval(reg_vprbs_tx_idi_driver_total_interval[15:0]),
				       .reg_vprbs_tx_idi_driver_virtual_channel(reg_vprbs_tx_idi_driver_virtual_channel[3:0]),
				       .reg_vprbs_tx_idi_driver_word_count(reg_vprbs_tx_idi_driver_word_count[15:0]),
				       .reg_vprbs_tx_mode(reg_vprbs_tx_mode[2:0]),
				       .reg_vprbs_tx_order(reg_vprbs_tx_order),
				       .reg_vprbs_tx_pat_reset(reg_vprbs_tx_pat_reset),
				       .idi_chk_header_en(as6s_csi_header_en), // Templated
				       .idi_chk_data_en	(as6s_csi_data_en), // Templated
				       .idi_chk_byte_en	(as6s_csi_bytes_en[2:0]), // Templated
				       .idi_chk_data_type(as6s_csi_data_type[5:0]), // Templated
				       .idi_chk_data	(as6s_csi_data[63:0]), // Templated
				       .reg_vprbs_loopback(reg_vprbs_loopback));





/*  vpg_idi  AUTO_TEMPLATE (
        .vpg_pkt_size_qst (vpg_pkt_size_qst@[]),
		.task_reg_vc_max(2'd0),
        .idi\(.*\)    (idi_vpg\1_lane@[]),
        .ppi\(.*\)    (ppi\10[]),
        .vpg\(.*\)    (vpg\1@[]),
		.ppi_clk      (ppi_clk@),
		.ppi_clkrstz  (ppi_clkrstz@),
)*/
vpg_idi u0_vpg_idi(/*autoinst*/
		   // Outputs
		   .idi_word_count	(idi_vpg_word_count_lane0[15:0]), // Templated
		   .idi_byte_en		(idi_vpg_byte_en_lane0[2:0]), // Templated
		   .idi_header_en	(idi_vpg_header_en_lane0), // Templated
		   .idi_data_en		(idi_vpg_data_en_lane0), // Templated
		   .idi_data		(idi_vpg_data_lane0[63:0]), // Templated
		   .idi_vc		(idi_vpg_vc_lane0[1:0]), // Templated
		   .idi_vcx		(idi_vpg_vcx_lane0[1:0]), // Templated
		   .idi_dt		(idi_vpg_dt_lane0[5:0]), // Templated
		   // Inputs
		   .ppi_clk		(ppi_clk0),		 // Templated
		   .ppi_clkrstz		(ppi_clkrstz0),		 // Templated
		   .vpg_bk_lines_qst	(vpg_bk_lines_qst0[`CSI2_DEVICE_VPG_BK_LINES_RS-1:0]), // Templated
		   .vpg_dt_qst		(vpg_dt_qst0[`CSI2_DEVICE_VPG_DT_RS-1:0]), // Templated
		   .vpg_en		(vpg_en0),		 // Templated
		   .vpg_frame_num_mode_qst(vpg_frame_num_mode_qst0[`CSI2_DEVICE_VPG_FRAME_NUM_MODE_RS-1:0]), // Templated
		   .vpg_hbp_time_qst	(vpg_hbp_time_qst0[`CSI2_DEVICE_VPG_HBP_TIME_RS-1:0]), // Templated
		   .vpg_hline_time_qst	(vpg_hline_time_qst0[`CSI2_DEVICE_VPG_HLINE_TIME_RS-1:0]), // Templated
		   .vpg_hsa_time_qst	(vpg_hsa_time_qst0[`CSI2_DEVICE_VPG_HSA_TIME_RS-1:0]), // Templated
		   .vpg_hsync_packet_en_qst(vpg_hsync_packet_en_qst0), // Templated
		   .vpg_line_num_mode_qst(vpg_line_num_mode_qst0[`CSI2_DEVICE_VPG_LINE_NUM_MODE_RS-1:0]), // Templated
		   .vpg_max_frame_num_qst(vpg_max_frame_num_qst0[`CSI2_DEVICE_VPG_MAX_FRAME_NUM_RS-1:0]), // Templated
		   .vpg_mode_qst	(vpg_mode_qst0),	 // Templated
		   .vpg_orientation_qst	(vpg_orientation_qst0),	 // Templated
		   .vpg_packet_lost_ack	(vpg_packet_lost_ack0),	 // Templated
		   .vpg_pkt_size_qst	(vpg_pkt_size_qst0[`CSI2_DEVICE_VPG_PKT_SIZE_RS-1:0]), // Templated
		   .vpg_start_line_num_qst(vpg_start_line_num_qst0[`CSI2_DEVICE_VPG_START_LINE_NUM_RS-1:0]), // Templated
		   .vpg_step_line_num_qst(vpg_step_line_num_qst0[`CSI2_DEVICE_VPG_STEP_LINE_NUM_RS-1:0]), // Templated
		   .vpg_vactive_lines_qst(vpg_vactive_lines_qst0[`CSI2_DEVICE_VPG_ACT_LINES_RS-1:0]), // Templated
		   .vpg_vbp_lines_qst	(vpg_vbp_lines_qst0[`CSI2_DEVICE_VPG_VBP_LINES_RS-1:0]), // Templated
		   .vpg_vc_qst		(vpg_vc_qst0[`CSI2_DEVICE_VPG_VC_RS-1:0]), // Templated
		   .vpg_vcx_qst		(vpg_vcx_qst0[`CSI2_DEVICE_VCX_DWIDTH-1:0]), // Templated
		   .vpg_vfp_lines_qst	(vpg_vfp_lines_qst0[`CSI2_DEVICE_VPG_VFP_LINES_RS-1:0]), // Templated
		   .vpg_vsa_lines_qst	(vpg_vsa_lines_qst0[`CSI2_DEVICE_VPG_VSA_LINES_RS-1:0]), // Templated
		   .task_reg_vc_max	(2'd0));			 // Templated

vpg_idi u1_vpg_idi(/*autoinst*/
		   // Outputs
		   .idi_word_count	(idi_vpg_word_count_lane1[15:0]), // Templated
		   .idi_byte_en		(idi_vpg_byte_en_lane1[2:0]), // Templated
		   .idi_header_en	(idi_vpg_header_en_lane1), // Templated
		   .idi_data_en		(idi_vpg_data_en_lane1), // Templated
		   .idi_data		(idi_vpg_data_lane1[63:0]), // Templated
		   .idi_vc		(idi_vpg_vc_lane1[1:0]), // Templated
		   .idi_vcx		(idi_vpg_vcx_lane1[1:0]), // Templated
		   .idi_dt		(idi_vpg_dt_lane1[5:0]), // Templated
		   // Inputs
		   .ppi_clk		(ppi_clk1),		 // Templated
		   .ppi_clkrstz		(ppi_clkrstz1),		 // Templated
		   .vpg_bk_lines_qst	(vpg_bk_lines_qst1[`CSI2_DEVICE_VPG_BK_LINES_RS-1:0]), // Templated
		   .vpg_dt_qst		(vpg_dt_qst1[`CSI2_DEVICE_VPG_DT_RS-1:0]), // Templated
		   .vpg_en		(vpg_en1),		 // Templated
		   .vpg_frame_num_mode_qst(vpg_frame_num_mode_qst1[`CSI2_DEVICE_VPG_FRAME_NUM_MODE_RS-1:0]), // Templated
		   .vpg_hbp_time_qst	(vpg_hbp_time_qst1[`CSI2_DEVICE_VPG_HBP_TIME_RS-1:0]), // Templated
		   .vpg_hline_time_qst	(vpg_hline_time_qst1[`CSI2_DEVICE_VPG_HLINE_TIME_RS-1:0]), // Templated
		   .vpg_hsa_time_qst	(vpg_hsa_time_qst1[`CSI2_DEVICE_VPG_HSA_TIME_RS-1:0]), // Templated
		   .vpg_hsync_packet_en_qst(vpg_hsync_packet_en_qst1), // Templated
		   .vpg_line_num_mode_qst(vpg_line_num_mode_qst1[`CSI2_DEVICE_VPG_LINE_NUM_MODE_RS-1:0]), // Templated
		   .vpg_max_frame_num_qst(vpg_max_frame_num_qst1[`CSI2_DEVICE_VPG_MAX_FRAME_NUM_RS-1:0]), // Templated
		   .vpg_mode_qst	(vpg_mode_qst1),	 // Templated
		   .vpg_orientation_qst	(vpg_orientation_qst1),	 // Templated
		   .vpg_packet_lost_ack	(vpg_packet_lost_ack1),	 // Templated
		   .vpg_pkt_size_qst	(vpg_pkt_size_qst1[`CSI2_DEVICE_VPG_PKT_SIZE_RS-1:0]), // Templated
		   .vpg_start_line_num_qst(vpg_start_line_num_qst1[`CSI2_DEVICE_VPG_START_LINE_NUM_RS-1:0]), // Templated
		   .vpg_step_line_num_qst(vpg_step_line_num_qst1[`CSI2_DEVICE_VPG_STEP_LINE_NUM_RS-1:0]), // Templated
		   .vpg_vactive_lines_qst(vpg_vactive_lines_qst1[`CSI2_DEVICE_VPG_ACT_LINES_RS-1:0]), // Templated
		   .vpg_vbp_lines_qst	(vpg_vbp_lines_qst1[`CSI2_DEVICE_VPG_VBP_LINES_RS-1:0]), // Templated
		   .vpg_vc_qst		(vpg_vc_qst1[`CSI2_DEVICE_VPG_VC_RS-1:0]), // Templated
		   .vpg_vcx_qst		(vpg_vcx_qst1[`CSI2_DEVICE_VCX_DWIDTH-1:0]), // Templated
		   .vpg_vfp_lines_qst	(vpg_vfp_lines_qst1[`CSI2_DEVICE_VPG_VFP_LINES_RS-1:0]), // Templated
		   .vpg_vsa_lines_qst	(vpg_vsa_lines_qst1[`CSI2_DEVICE_VPG_VSA_LINES_RS-1:0]), // Templated
		   .task_reg_vc_max	(2'd0));			 // Templated

vpg_idi u2_vpg_idi(/*autoinst*/
		   // Outputs
		   .idi_word_count	(idi_vpg_word_count_lane2[15:0]), // Templated
		   .idi_byte_en		(idi_vpg_byte_en_lane2[2:0]), // Templated
		   .idi_header_en	(idi_vpg_header_en_lane2), // Templated
		   .idi_data_en		(idi_vpg_data_en_lane2), // Templated
		   .idi_data		(idi_vpg_data_lane2[63:0]), // Templated
		   .idi_vc		(idi_vpg_vc_lane2[1:0]), // Templated
		   .idi_vcx		(idi_vpg_vcx_lane2[1:0]), // Templated
		   .idi_dt		(idi_vpg_dt_lane2[5:0]), // Templated
		   // Inputs
		   .ppi_clk		(ppi_clk2),		 // Templated
		   .ppi_clkrstz		(ppi_clkrstz2),		 // Templated
		   .vpg_bk_lines_qst	(vpg_bk_lines_qst2[`CSI2_DEVICE_VPG_BK_LINES_RS-1:0]), // Templated
		   .vpg_dt_qst		(vpg_dt_qst2[`CSI2_DEVICE_VPG_DT_RS-1:0]), // Templated
		   .vpg_en		(vpg_en2),		 // Templated
		   .vpg_frame_num_mode_qst(vpg_frame_num_mode_qst2[`CSI2_DEVICE_VPG_FRAME_NUM_MODE_RS-1:0]), // Templated
		   .vpg_hbp_time_qst	(vpg_hbp_time_qst2[`CSI2_DEVICE_VPG_HBP_TIME_RS-1:0]), // Templated
		   .vpg_hline_time_qst	(vpg_hline_time_qst2[`CSI2_DEVICE_VPG_HLINE_TIME_RS-1:0]), // Templated
		   .vpg_hsa_time_qst	(vpg_hsa_time_qst2[`CSI2_DEVICE_VPG_HSA_TIME_RS-1:0]), // Templated
		   .vpg_hsync_packet_en_qst(vpg_hsync_packet_en_qst2), // Templated
		   .vpg_line_num_mode_qst(vpg_line_num_mode_qst2[`CSI2_DEVICE_VPG_LINE_NUM_MODE_RS-1:0]), // Templated
		   .vpg_max_frame_num_qst(vpg_max_frame_num_qst2[`CSI2_DEVICE_VPG_MAX_FRAME_NUM_RS-1:0]), // Templated
		   .vpg_mode_qst	(vpg_mode_qst2),	 // Templated
		   .vpg_orientation_qst	(vpg_orientation_qst2),	 // Templated
		   .vpg_packet_lost_ack	(vpg_packet_lost_ack2),	 // Templated
		   .vpg_pkt_size_qst	(vpg_pkt_size_qst2[`CSI2_DEVICE_VPG_PKT_SIZE_RS-1:0]), // Templated
		   .vpg_start_line_num_qst(vpg_start_line_num_qst2[`CSI2_DEVICE_VPG_START_LINE_NUM_RS-1:0]), // Templated
		   .vpg_step_line_num_qst(vpg_step_line_num_qst2[`CSI2_DEVICE_VPG_STEP_LINE_NUM_RS-1:0]), // Templated
		   .vpg_vactive_lines_qst(vpg_vactive_lines_qst2[`CSI2_DEVICE_VPG_ACT_LINES_RS-1:0]), // Templated
		   .vpg_vbp_lines_qst	(vpg_vbp_lines_qst2[`CSI2_DEVICE_VPG_VBP_LINES_RS-1:0]), // Templated
		   .vpg_vc_qst		(vpg_vc_qst2[`CSI2_DEVICE_VPG_VC_RS-1:0]), // Templated
		   .vpg_vcx_qst		(vpg_vcx_qst2[`CSI2_DEVICE_VCX_DWIDTH-1:0]), // Templated
		   .vpg_vfp_lines_qst	(vpg_vfp_lines_qst2[`CSI2_DEVICE_VPG_VFP_LINES_RS-1:0]), // Templated
		   .vpg_vsa_lines_qst	(vpg_vsa_lines_qst2[`CSI2_DEVICE_VPG_VSA_LINES_RS-1:0]), // Templated
		   .task_reg_vc_max	(2'd0));			 // Templated

vpg_idi u3_vpg_idi(/*autoinst*/
		   // Outputs
		   .idi_word_count	(idi_vpg_word_count_lane3[15:0]), // Templated
		   .idi_byte_en		(idi_vpg_byte_en_lane3[2:0]), // Templated
		   .idi_header_en	(idi_vpg_header_en_lane3), // Templated
		   .idi_data_en		(idi_vpg_data_en_lane3), // Templated
		   .idi_data		(idi_vpg_data_lane3[63:0]), // Templated
		   .idi_vc		(idi_vpg_vc_lane3[1:0]), // Templated
		   .idi_vcx		(idi_vpg_vcx_lane3[1:0]), // Templated
		   .idi_dt		(idi_vpg_dt_lane3[5:0]), // Templated
		   // Inputs
		   .ppi_clk		(ppi_clk3),		 // Templated
		   .ppi_clkrstz		(ppi_clkrstz3),		 // Templated
		   .vpg_bk_lines_qst	(vpg_bk_lines_qst3[`CSI2_DEVICE_VPG_BK_LINES_RS-1:0]), // Templated
		   .vpg_dt_qst		(vpg_dt_qst3[`CSI2_DEVICE_VPG_DT_RS-1:0]), // Templated
		   .vpg_en		(vpg_en3),		 // Templated
		   .vpg_frame_num_mode_qst(vpg_frame_num_mode_qst3[`CSI2_DEVICE_VPG_FRAME_NUM_MODE_RS-1:0]), // Templated
		   .vpg_hbp_time_qst	(vpg_hbp_time_qst3[`CSI2_DEVICE_VPG_HBP_TIME_RS-1:0]), // Templated
		   .vpg_hline_time_qst	(vpg_hline_time_qst3[`CSI2_DEVICE_VPG_HLINE_TIME_RS-1:0]), // Templated
		   .vpg_hsa_time_qst	(vpg_hsa_time_qst3[`CSI2_DEVICE_VPG_HSA_TIME_RS-1:0]), // Templated
		   .vpg_hsync_packet_en_qst(vpg_hsync_packet_en_qst3), // Templated
		   .vpg_line_num_mode_qst(vpg_line_num_mode_qst3[`CSI2_DEVICE_VPG_LINE_NUM_MODE_RS-1:0]), // Templated
		   .vpg_max_frame_num_qst(vpg_max_frame_num_qst3[`CSI2_DEVICE_VPG_MAX_FRAME_NUM_RS-1:0]), // Templated
		   .vpg_mode_qst	(vpg_mode_qst3),	 // Templated
		   .vpg_orientation_qst	(vpg_orientation_qst3),	 // Templated
		   .vpg_packet_lost_ack	(vpg_packet_lost_ack3),	 // Templated
		   .vpg_pkt_size_qst	(vpg_pkt_size_qst3[`CSI2_DEVICE_VPG_PKT_SIZE_RS-1:0]), // Templated
		   .vpg_start_line_num_qst(vpg_start_line_num_qst3[`CSI2_DEVICE_VPG_START_LINE_NUM_RS-1:0]), // Templated
		   .vpg_step_line_num_qst(vpg_step_line_num_qst3[`CSI2_DEVICE_VPG_STEP_LINE_NUM_RS-1:0]), // Templated
		   .vpg_vactive_lines_qst(vpg_vactive_lines_qst3[`CSI2_DEVICE_VPG_ACT_LINES_RS-1:0]), // Templated
		   .vpg_vbp_lines_qst	(vpg_vbp_lines_qst3[`CSI2_DEVICE_VPG_VBP_LINES_RS-1:0]), // Templated
		   .vpg_vc_qst		(vpg_vc_qst3[`CSI2_DEVICE_VPG_VC_RS-1:0]), // Templated
		   .vpg_vcx_qst		(vpg_vcx_qst3[`CSI2_DEVICE_VCX_DWIDTH-1:0]), // Templated
		   .vpg_vfp_lines_qst	(vpg_vfp_lines_qst3[`CSI2_DEVICE_VPG_VFP_LINES_RS-1:0]), // Templated
		   .vpg_vsa_lines_qst	(vpg_vsa_lines_qst3[`CSI2_DEVICE_VPG_VSA_LINES_RS-1:0]), // Templated
		   .task_reg_vc_max	(2'd0));			 // Templated


wire [3:0]                        cnt_line_end_rd_side0             ;
wire [3:0]                        cnt_line_end_rd_side1             ;    
wire [3:0]                        cnt_line_end_rd_side2             ;    
wire [3:0]                        cnt_line_end_rd_side3             ;    
wire [2:0]                        fifo_rd_ctrl_cs0                  ;   
wire [2:0]                        fifo_rd_ctrl_cs1                  ;   
wire [2:0]                        fifo_rd_ctrl_cs2                  ;   
wire [2:0]                        fifo_rd_ctrl_cs3                  ;   
wire                            fs_detect_pipe0                     ;    
wire                            fs_detect_pipe1                     ;    
wire                            fs_detect_pipe2                     ;    
wire                            fs_detect_pipe3                     ;    
wire [1:0]        to_clkgen_fifo_rdclk_sel0;// From u0_as6d_app_fifo_rdclk_sel of as6d_app_fifo_rdclk_sel.v
wire [1:0]        to_clkgen_fifo_rdclk_sel1;// From u1_as6d_app_fifo_rdclk_sel of as6d_app_fifo_rdclk_sel.v
wire [1:0]        to_clkgen_fifo_rdclk_sel2;// From u2_as6d_app_fifo_rdclk_sel of as6d_app_fifo_rdclk_sel.v
wire [1:0]        to_clkgen_fifo_rdclk_sel3;// From u3_as6d_app_fifo_rdclk_sel of as6d_app_fifo_rdclk_sel.v
wire    [1:0]        to_clkgen_fifo_wrclk_sel0    ;
wire    [1:0]        to_clkgen_fifo_wrclk_sel1    ;
wire    [1:0]        to_clkgen_fifo_wrclk_sel2    ;
wire    [1:0]        to_clkgen_fifo_wrclk_sel3    ;
wire [9:0]        reg_dft_sync_tpram_config;// To u_as6d_app_video_pipe of as6d_app_video_pipe.v
wire [8:0]        reg_dft_tpram_config;    // To u_as6d_app_video_pipe of as6d_app_video_pipe.v
wire            reg_testbus_hi8bsel_8bmode;// To u_as6d_app_mon_top of as6d_app_mon_top.v
wire [15:0]                        reg_rd_dig_test_bus;    // From u_as6d_app_mon_top of as6d_app_mon_top.v
wire [5:0]        reg_testbus_sel_hi0;    // To u_as6d_app_mon_top of as6d_app_mon_top.v
wire [5:0]        reg_testbus_sel_hi1;    // To u_as6d_app_mon_top of as6d_app_mon_top.v
wire [5:0]        reg_testbus_sel_lo0;    // To u_as6d_app_mon_top of as6d_app_mon_top.v
wire [5:0]        reg_testbus_sel_lo1;    // To u_as6d_app_mon_top of as6d_app_mon_top.v
wire [3:0]        reg_testbus_sel_order0;    // To u_as6d_app_mon_top of as6d_app_mon_top.v
wire [3:0]        reg_testbus_sel_order1;    // To u_as6d_app_mon_top of as6d_app_mon_top.v
wire [15:0]        reg_testbus_sel_swap;    // To u_as6d_app_mon_top of as6d_app_mon_top.v
wire [15:0]        PIN_DIG_TEST_BUS;    // From u_as6d_app_mon_top of as6d_app_mon_top.v

/*as6d_app    AUTO_TEMPLATE(
        .mep\(.*\)_byte_en              (idi_byte_en_lane\1[]),
        .mep\(.*\)_csi_data             (idi_data_lane\1[]),
        .mep\(.*\)_data_en              (idi_data_en_lane\1),
        .mep\(.*\)_data_type            (idi_dt_lane\1[]),
        .mep\(.*\)_header_en            (idi_header_en_lane\1),
        .mep\(.*\)_virtual_channel      (idi_vc_lane\1[]),
        .mep\(.*\)_virtual_channel_x    (idi_vcx_lane\1[]),
        .mep\(.*\)_word_count           (idi_word_count_lane\1[]),
		.mep\(.*\)_tunnel_mode_en       (1'd0),


        .reg_pipe1_map_en               (reg_pipe1_map_en),

		.aggr0_idi_\(.*\)(idi_prbs_chk_\1[]),

        .to_clkgen_fifo_rdclk_sel\(.*\)    (),
        .to_clkgen_fifo_wrclk_sel\(.*\)    (),
        .aggr\(.*\)_idi\(.*\)                    (),
        .reg_pipe0_map0_aggr_id    (reg_pipe0_map0_aggr_id),
        .reg_pipe0_map1_aggr_id    (reg_pipe0_map1_aggr_id),
        .reg_pipe0_map2_aggr_id    (reg_pipe0_map2_aggr_id),
        .reg_pipe0_map3_aggr_id    (reg_pipe0_map3_aggr_id),
        .reg_pipe0_map4_aggr_id    (reg_pipe0_map4_aggr_id),
        .reg_pipe0_map5_aggr_id    (reg_pipe0_map5_aggr_id),
        .reg_pipe0_map6_aggr_id    (reg_pipe0_map6_aggr_id),
        .reg_pipe0_map7_aggr_id    (reg_pipe0_map7_aggr_id),
        .reg_pipe0_map8_aggr_id    (reg_pipe0_map8_aggr_id),
        .reg_pipe0_map9_aggr_id    (reg_pipe0_map9_aggr_id),
        .reg_pipe0_map10_aggr_id(reg_pipe0_map10_aggr_id),
        .reg_pipe0_map11_aggr_id(reg_pipe0_map11_aggr_id),
        .reg_pipe0_map12_aggr_id(reg_pipe0_map12_aggr_id),
        .reg_pipe0_map13_aggr_id(reg_pipe0_map13_aggr_id),
        .reg_pipe0_map14_aggr_id(reg_pipe0_map14_aggr_id),
        .reg_pipe0_map15_aggr_id(reg_pipe0_map15_aggr_id),
        .reg_pipe1_map0_aggr_id    (reg_pipe1_map0_aggr_id),
        .reg_pipe1_map1_aggr_id    (reg_pipe1_map1_aggr_id),
        .reg_pipe1_map2_aggr_id    (reg_pipe1_map2_aggr_id),
        .reg_pipe1_map3_aggr_id    (reg_pipe1_map3_aggr_id),
        .reg_pipe1_map4_aggr_id    (reg_pipe1_map4_aggr_id),
        .reg_pipe1_map5_aggr_id    (reg_pipe1_map5_aggr_id),
        .reg_pipe1_map6_aggr_id    (reg_pipe1_map6_aggr_id),
        .reg_pipe1_map7_aggr_id    (reg_pipe1_map7_aggr_id),
        .reg_pipe1_map8_aggr_id    (reg_pipe1_map8_aggr_id),
        .reg_pipe1_map9_aggr_id    (reg_pipe1_map9_aggr_id),
        .reg_pipe1_map10_aggr_id(reg_pipe1_map10_aggr_id),
        .reg_pipe1_map11_aggr_id(reg_pipe1_map11_aggr_id),
        .reg_pipe1_map12_aggr_id(reg_pipe1_map12_aggr_id),
        .reg_pipe1_map13_aggr_id(reg_pipe1_map13_aggr_id),
        .reg_pipe1_map14_aggr_id(reg_pipe1_map14_aggr_id),
        .reg_pipe1_map15_aggr_id(reg_pipe1_map15_aggr_id),
        .reg_pipe2_map0_aggr_id    (reg_pipe2_map0_aggr_id),
        .reg_pipe2_map1_aggr_id    (reg_pipe2_map1_aggr_id),
        .reg_pipe2_map2_aggr_id    (reg_pipe2_map2_aggr_id),
        .reg_pipe2_map3_aggr_id    (reg_pipe2_map3_aggr_id),
        .reg_pipe2_map4_aggr_id    (reg_pipe2_map4_aggr_id),
        .reg_pipe2_map5_aggr_id    (reg_pipe2_map5_aggr_id),
        .reg_pipe2_map6_aggr_id    (reg_pipe2_map6_aggr_id),
        .reg_pipe2_map7_aggr_id    (reg_pipe2_map7_aggr_id),
        .reg_pipe2_map8_aggr_id    (reg_pipe2_map8_aggr_id),
        .reg_pipe2_map9_aggr_id    (reg_pipe2_map9_aggr_id),
        .reg_pipe2_map10_aggr_id(reg_pipe2_map10_aggr_id),
        .reg_pipe2_map11_aggr_id(reg_pipe2_map11_aggr_id),
        .reg_pipe2_map12_aggr_id(reg_pipe2_map12_aggr_id),
        .reg_pipe2_map13_aggr_id(reg_pipe2_map13_aggr_id),
        .reg_pipe2_map14_aggr_id(reg_pipe2_map14_aggr_id),
        .reg_pipe2_map15_aggr_id(reg_pipe2_map15_aggr_id),
        .reg_pipe3_map0_aggr_id    (reg_pipe3_map0_aggr_id),
        .reg_pipe3_map1_aggr_id    (reg_pipe3_map1_aggr_id),
        .reg_pipe3_map2_aggr_id    (reg_pipe3_map2_aggr_id),
        .reg_pipe3_map3_aggr_id    (reg_pipe3_map3_aggr_id),
        .reg_pipe3_map4_aggr_id    (reg_pipe3_map4_aggr_id),
        .reg_pipe3_map5_aggr_id    (reg_pipe3_map5_aggr_id),
        .reg_pipe3_map6_aggr_id    (reg_pipe3_map6_aggr_id),
        .reg_pipe3_map7_aggr_id    (reg_pipe3_map7_aggr_id),
        .reg_pipe3_map8_aggr_id    (reg_pipe3_map8_aggr_id),
        .reg_pipe3_map9_aggr_id    (reg_pipe3_map9_aggr_id),
        .reg_pipe3_map10_aggr_id(reg_pipe3_map10_aggr_id),
        .reg_pipe3_map11_aggr_id(reg_pipe3_map11_aggr_id),
        .reg_pipe3_map12_aggr_id(reg_pipe3_map12_aggr_id),
        .reg_pipe3_map13_aggr_id(reg_pipe3_map13_aggr_id),
        .reg_pipe3_map14_aggr_id(reg_pipe3_map14_aggr_id),
        .reg_pipe3_map15_aggr_id(reg_pipe3_map15_aggr_id),
        .reg_pipe\(.*\)_map0_vc_source (reg_pipe\1_map0_vc_source ),            
        .reg_pipe\(.*\)_map1_vc_source (reg_pipe\1_map1_vc_source ),            
        .reg_pipe\(.*\)_map2_vc_source (reg_pipe\1_map2_vc_source ),            
        .reg_pipe\(.*\)_map3_vc_source (reg_pipe\1_map3_vc_source ),            
        .reg_pipe\(.*\)_map4_vc_source (reg_pipe\1_map4_vc_source ),            
        .reg_pipe\(.*\)_map5_vc_source (reg_pipe\1_map5_vc_source ),            
        .reg_pipe\(.*\)_map6_vc_source (reg_pipe\1_map6_vc_source ),            
        .reg_pipe\(.*\)_map7_vc_source (reg_pipe\1_map7_vc_source ),            
        .reg_pipe\(.*\)_map8_vc_source (reg_pipe\1_map8_vc_source ),            
        .reg_pipe\(.*\)_map9_vc_source (reg_pipe\1_map9_vc_source ),            
        .reg_pipe\(.*\)_map10_vc_source(reg_pipe\1_map10_vc_source),            
        .reg_pipe\(.*\)_map11_vc_source(reg_pipe\1_map11_vc_source),            
        .reg_pipe\(.*\)_map12_vc_source(reg_pipe\1_map12_vc_source),            
        .reg_pipe\(.*\)_map13_vc_source(reg_pipe\1_map13_vc_source),            
        .reg_pipe\(.*\)_map14_vc_source(reg_pipe\1_map14_vc_source),            
        .reg_pipe\(.*\)_map15_vc_source(reg_pipe\1_map15_vc_source),            
        .reg_pipe\(.*\)_map0_vc_dest (reg_pipe\1_map0_vc_dest )      ,      
        .reg_pipe\(.*\)_map1_vc_dest (reg_pipe\1_map1_vc_dest )      ,      
        .reg_pipe\(.*\)_map2_vc_dest (reg_pipe\1_map2_vc_dest )      ,      
        .reg_pipe\(.*\)_map3_vc_dest (reg_pipe\1_map3_vc_dest )      ,      
        .reg_pipe\(.*\)_map4_vc_dest (reg_pipe\1_map4_vc_dest )      ,      
        .reg_pipe\(.*\)_map5_vc_dest (reg_pipe\1_map5_vc_dest )      ,      
        .reg_pipe\(.*\)_map6_vc_dest (reg_pipe\1_map6_vc_dest )      ,      
        .reg_pipe\(.*\)_map7_vc_dest (reg_pipe\1_map7_vc_dest )      ,      
        .reg_pipe\(.*\)_map8_vc_dest (reg_pipe\1_map8_vc_dest )      ,      
        .reg_pipe\(.*\)_map9_vc_dest (reg_pipe\1_map9_vc_dest )      ,      
        .reg_pipe\(.*\)_map10_vc_dest(reg_pipe\1_map10_vc_dest)      ,      
        .reg_pipe\(.*\)_map11_vc_dest(reg_pipe\1_map11_vc_dest)      ,      
        .reg_pipe\(.*\)_map12_vc_dest(reg_pipe\1_map12_vc_dest)      ,      
        .reg_pipe\(.*\)_map13_vc_dest(reg_pipe\1_map13_vc_dest)      ,      
        .reg_pipe\(.*\)_map14_vc_dest(reg_pipe\1_map14_vc_dest)      ,      
        .reg_pipe\(.*\)_map15_vc_dest(reg_pipe\1_map15_vc_dest)      ,      
        .reg_pipe\(.*\)_map0_dt_source (reg_pipe\1_map0_dt_source ),            
        .reg_pipe\(.*\)_map1_dt_source (reg_pipe\1_map1_dt_source ),            
        .reg_pipe\(.*\)_map2_dt_source (reg_pipe\1_map2_dt_source ),            
        .reg_pipe\(.*\)_map3_dt_source (reg_pipe\1_map3_dt_source ),            
        .reg_pipe\(.*\)_map4_dt_source (reg_pipe\1_map4_dt_source ),            
        .reg_pipe\(.*\)_map5_dt_source (reg_pipe\1_map5_dt_source ),            
        .reg_pipe\(.*\)_map6_dt_source (reg_pipe\1_map6_dt_source ),            
        .reg_pipe\(.*\)_map7_dt_source (reg_pipe\1_map7_dt_source ),            
        .reg_pipe\(.*\)_map8_dt_source (reg_pipe\1_map8_dt_source ),            
        .reg_pipe\(.*\)_map9_dt_source (reg_pipe\1_map9_dt_source ),            
        .reg_pipe\(.*\)_map10_dt_source(reg_pipe\1_map10_dt_source),            
        .reg_pipe\(.*\)_map11_dt_source(reg_pipe\1_map11_dt_source),            
        .reg_pipe\(.*\)_map12_dt_source(reg_pipe\1_map12_dt_source),            
        .reg_pipe\(.*\)_map13_dt_source(reg_pipe\1_map13_dt_source),            
        .reg_pipe\(.*\)_map14_dt_source(reg_pipe\1_map14_dt_source),            
        .reg_pipe\(.*\)_map15_dt_source(reg_pipe\1_map15_dt_source),            
        .reg_pipe\(.*\)_map0_dt_dest (reg_pipe\1_map0_dt_dest ),            
        .reg_pipe\(.*\)_map1_dt_dest (reg_pipe\1_map1_dt_dest ),            
        .reg_pipe\(.*\)_map2_dt_dest (reg_pipe\1_map2_dt_dest ),            
        .reg_pipe\(.*\)_map3_dt_dest (reg_pipe\1_map3_dt_dest ),            
        .reg_pipe\(.*\)_map4_dt_dest (reg_pipe\1_map4_dt_dest ),            
        .reg_pipe\(.*\)_map5_dt_dest (reg_pipe\1_map5_dt_dest ),            
        .reg_pipe\(.*\)_map6_dt_dest (reg_pipe\1_map6_dt_dest ),            
        .reg_pipe\(.*\)_map7_dt_dest (reg_pipe\1_map7_dt_dest ),            
        .reg_pipe\(.*\)_map8_dt_dest (reg_pipe\1_map8_dt_dest ),            
        .reg_pipe\(.*\)_map9_dt_dest (reg_pipe\1_map9_dt_dest ),            
        .reg_pipe\(.*\)_map10_dt_dest(reg_pipe\1_map10_dt_dest),            
        .reg_pipe\(.*\)_map11_dt_dest(reg_pipe\1_map11_dt_dest),            
        .reg_pipe\(.*\)_map12_dt_dest(reg_pipe\1_map12_dt_dest),            
        .reg_pipe\(.*\)_map13_dt_dest(reg_pipe\1_map13_dt_dest),            
        .reg_pipe\(.*\)_map14_dt_dest(reg_pipe\1_map14_dt_dest),            
        .reg_pipe\(.*\)_map15_dt_dest(reg_pipe\1_map15_dt_dest),            
        .reg_pipe\(.*\)_map_en            (reg_pipe\1_map_en),
        .reg_rd_fifo_rd_ctrl_cs\(.*\)(),
        .reg_rd_fs_cnt_pipe\(.*\)    (),
        .reg_rd_cnt_line_end_rd_side\(.*\)(),
        .reg_rd_sch0_cs    (),
        .reg_rd_sch1_cs    (),
        .reg_rd_sch2_cs    (),
        .reg_rd_sch3_cs    (),

        .reg_resv_pkt_match_lp_dt_en\(.*\)   (reg_resv_pkt_match_lp_dt_en ),
        .reg_resv_pkt_match_lp_dt\(.*\)      (reg_resv_pkt_match_lp_dt    ),
        .reg_clear_resv_pkt_cnt_lp_pf\(.*\)  (reg_clear_resv_pkt_cnt_lp_pf),
        .reg_clear_resv_pkt_cnt_lp_ph\(.*\)  (reg_clear_resv_pkt_cnt_lp_ph),
        .reg_clear_resv_pkt_cnt_sp_fe\(.*\)  (reg_clear_resv_pkt_cnt_sp_fe),
        .reg_clear_resv_pkt_cnt_sp_fs\(.*\)  (reg_clear_resv_pkt_cnt_sp_fs),
        .reg_clear_resv_pkt_cnt_sp_le\(.*\)  (reg_clear_resv_pkt_cnt_sp_le),
        .reg_clear_resv_pkt_cnt_sp_ls\(.*\)  (reg_clear_resv_pkt_cnt_sp_ls),
        .reg_send_pkt_match_lp_dt_en\(.*\)   (reg_send_pkt_match_lp_dt_en ),
        .reg_send_pkt_match_lp_dt\(.*\)      (reg_send_pkt_match_lp_dt    ),
        .reg_clear_send_pkt_cnt_lp_pf\(.*\)  (reg_clear_send_pkt_cnt_lp_pf),
        .reg_clear_send_pkt_cnt_lp_ph\(.*\)  (reg_clear_send_pkt_cnt_lp_ph),
        .reg_clear_send_pkt_cnt_sp_fe\(.*\)  (reg_clear_send_pkt_cnt_sp_fe),
        .reg_clear_send_pkt_cnt_sp_fs\(.*\)  (reg_clear_send_pkt_cnt_sp_fs),
        .reg_clear_send_pkt_cnt_sp_le\(.*\)  (reg_clear_send_pkt_cnt_sp_le),
        .reg_clear_send_pkt_cnt_sp_ls\(.*\)  (reg_clear_send_pkt_cnt_sp_ls),

        .reg_rd_resv_pkt_cnt\(.*\)  (),
        .reg_rd_send_pkt_cnt\(.*\)  (),

        .reg_rd_vprbs_rx_\(.*\)	(),
        .reg_vprbs_\(.*\)_app_route_lane\(.*\)	(reg_vprbs_\1[]),

		.reg_mem_dt\(.*\)_selz_mep\(.*\)	(reg_mem_dt\1_selz[]),
		.reg_mem_dt\(.*\)_selz_en_mep\(.*\)   (reg_mem_dt\1_selz_en),
		.reg_vc_selz_l_mep\(.*\)	(reg_vc_selz_l[]),
		.reg_vc_selz_h_mep\(.*\)	(reg_vc_selz_h[]),
        .mep_clk_rst_n\(.*\) (ppi_clkrstz\1),
        .mep_clk\(.*\) (ppi_clk\1),
		.reg_mep\(.*\)_tdi_en	(1'd0),
		.reg_mep\(.*\)_tdi_en_force(1'd0),
		.reg_dft_sync_tpram_config(10'd0),
		.reg_dft_tpram_config(9'd0),
		.reg_app_ecc_addr_protect_en(1'd1),
		.reg_app_ecc_bypass(1'd0),
		.reg_app_ecc_fault_detc_en(1'd1),
		.app_aggr_idi_crc_err_int0(),
		.app_aggr_idi_crc_err_int1(),
		.app_aggr_idi_crc_err_int2(),
		.app_aggr_idi_crc_err_int3(),
		.vprbs_rx_fail_app_route_int0(),
		.vprbs_rx_fail_app_route_int1(),
		.vprbs_rx_fail_app_route_int2(),
		.vprbs_rx_fail_app_route_int3(),
		.vprbs_rx_fail_app_route_int4(),
		.vprbs_rx_fail_app_route_int5(),
		.vprbs_rx_fail_app_route_int6(),
		.vprbs_rx_fail_app_route_int7(),
		.video_data_afifo_ovf_int0(video_data_afifo_ovf_int0),
		.video_data_afifo_ovf_int1(video_data_afifo_ovf_int1),
		.video_data_afifo_ovf_int2(video_data_afifo_ovf_int2),
		.video_data_afifo_ovf_int3(video_data_afifo_ovf_int3),
		.video_data_afifo_ovf_int4(video_data_afifo_ovf_int4),
		.video_data_afifo_ovf_int5(video_data_afifo_ovf_int5),
		.video_data_afifo_ovf_int6(video_data_afifo_ovf_int6),
		.video_data_afifo_ovf_int7(video_data_afifo_ovf_int7),
		.reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold(16'd200),
		.reg_dbg_pkt_num_nonzero_threshold(16'd200),
		.reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err(),
		.reg_rd_dbg_pkt_num_nonzero_threshold_err(),
		.reg_dbg_fcfs_method_2_mechine_en(1'd1),
		.reg_sch_data_type_align_fail_int_mask0(1'd0),
		.reg_sch_data_type_align_fail_int_mask1(1'd0),
		.reg_sch_data_type_align_fail_int_mask2(1'd0),
		.reg_sch_data_type_align_fail_int_mask3(1'd0),
);*/
as6d_app    u_as6d_app(/*AUTOINST*/
		       // Outputs
		       .PIN_DIG_TEST_BUS(PIN_DIG_TEST_BUS[15:0]),
		       .aggr0_idi_byte_en(idi_prbs_chk_byte_en[3:0]), // Templated
		       .aggr0_idi_data	(idi_prbs_chk_data[`CSI2_DEVICE_IDI_DATA_WIDTH-1:0]), // Templated
		       .aggr0_idi_data_en(idi_prbs_chk_data_en), // Templated
		       .aggr0_idi_data_parity(idi_prbs_chk_data_parity[20:0]), // Templated
		       .aggr0_idi_data_type(idi_prbs_chk_data_type[5:0]), // Templated
		       .aggr0_idi_header_en(idi_prbs_chk_header_en), // Templated
		       .aggr0_idi_tunnel_mode_en(idi_prbs_chk_tunnel_mode_en), // Templated
		       .aggr0_idi_virtual_channel(idi_prbs_chk_virtual_channel[1:0]), // Templated
		       .aggr0_idi_virtual_channel_x(idi_prbs_chk_virtual_channel_x[`CSI2_DEVICE_VCX_DWIDTH-1:0]), // Templated
		       .aggr0_idi_word_count(idi_prbs_chk_word_count[15:0]), // Templated
		       .aggr1_idi_byte_en(),			 // Templated
		       .aggr1_idi_data	(),			 // Templated
		       .aggr1_idi_data_en(),			 // Templated
		       .aggr1_idi_data_parity(),		 // Templated
		       .aggr1_idi_data_type(),			 // Templated
		       .aggr1_idi_header_en(),			 // Templated
		       .aggr1_idi_tunnel_mode_en(),		 // Templated
		       .aggr1_idi_virtual_channel(),		 // Templated
		       .aggr1_idi_virtual_channel_x(),		 // Templated
		       .aggr1_idi_word_count(),			 // Templated
		       .aggr2_idi_byte_en(),			 // Templated
		       .aggr2_idi_data	(),			 // Templated
		       .aggr2_idi_data_en(),			 // Templated
		       .aggr2_idi_data_parity(),		 // Templated
		       .aggr2_idi_data_type(),			 // Templated
		       .aggr2_idi_header_en(),			 // Templated
		       .aggr2_idi_tunnel_mode_en(),		 // Templated
		       .aggr2_idi_virtual_channel(),		 // Templated
		       .aggr2_idi_virtual_channel_x(),		 // Templated
		       .aggr2_idi_word_count(),			 // Templated
		       .aggr3_idi_byte_en(),			 // Templated
		       .aggr3_idi_data	(),			 // Templated
		       .aggr3_idi_data_en(),			 // Templated
		       .aggr3_idi_data_parity(),		 // Templated
		       .aggr3_idi_data_type(),			 // Templated
		       .aggr3_idi_header_en(),			 // Templated
		       .aggr3_idi_tunnel_mode_en(),		 // Templated
		       .aggr3_idi_virtual_channel(),		 // Templated
		       .aggr3_idi_virtual_channel_x(),		 // Templated
		       .aggr3_idi_word_count(),			 // Templated
		       .app_aggr_idi_crc_err_int0(),		 // Templated
		       .app_aggr_idi_crc_err_int1(),		 // Templated
		       .app_aggr_idi_crc_err_int2(),		 // Templated
		       .app_aggr_idi_crc_err_int3(),		 // Templated
		       .app_async_rst_req(app_async_rst_req),
		       .reg_rd_app_full_cnt_async_fifo_pipe0(reg_rd_app_full_cnt_async_fifo_pipe0[31:0]),
		       .reg_rd_app_full_cnt_async_fifo_pipe1(reg_rd_app_full_cnt_async_fifo_pipe1[31:0]),
		       .reg_rd_app_full_cnt_async_fifo_pipe2(reg_rd_app_full_cnt_async_fifo_pipe2[31:0]),
		       .reg_rd_app_full_cnt_async_fifo_pipe3(reg_rd_app_full_cnt_async_fifo_pipe3[31:0]),
		       .reg_rd_app_full_cnt_async_fifo_pipe4(reg_rd_app_full_cnt_async_fifo_pipe4[31:0]),
		       .reg_rd_app_full_cnt_async_fifo_pipe5(reg_rd_app_full_cnt_async_fifo_pipe5[31:0]),
		       .reg_rd_app_full_cnt_async_fifo_pipe6(reg_rd_app_full_cnt_async_fifo_pipe6[31:0]),
		       .reg_rd_app_full_cnt_async_fifo_pipe7(reg_rd_app_full_cnt_async_fifo_pipe7[31:0]),
		       .reg_rd_app_full_cnt_sync_fifo_pipe0(reg_rd_app_full_cnt_sync_fifo_pipe0[31:0]),
		       .reg_rd_app_full_cnt_sync_fifo_pipe1(reg_rd_app_full_cnt_sync_fifo_pipe1[31:0]),
		       .reg_rd_app_full_cnt_sync_fifo_pipe2(reg_rd_app_full_cnt_sync_fifo_pipe2[31:0]),
		       .reg_rd_app_full_cnt_sync_fifo_pipe3(reg_rd_app_full_cnt_sync_fifo_pipe3[31:0]),
		       .reg_rd_app_full_cnt_sync_fifo_pipe4(reg_rd_app_full_cnt_sync_fifo_pipe4[31:0]),
		       .reg_rd_app_full_cnt_sync_fifo_pipe5(reg_rd_app_full_cnt_sync_fifo_pipe5[31:0]),
		       .reg_rd_app_full_cnt_sync_fifo_pipe6(reg_rd_app_full_cnt_sync_fifo_pipe6[31:0]),
		       .reg_rd_app_full_cnt_sync_fifo_pipe7(reg_rd_app_full_cnt_sync_fifo_pipe7[31:0]),
		       .reg_rd_dbg_pkt_num_nonzero_and_fifo_empty_threshold_err(), // Templated
		       .reg_rd_dbg_pkt_num_nonzero_threshold_err(), // Templated
		       .reg_rd_dig_test_bus(reg_rd_dig_test_bus[15:0]),
		       .reg_rd_pipe_fifo_full(reg_rd_pipe_fifo_full[7:0]),
		       .reg_rd_resv_pkt_cnt_lp_pf_pipe0(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_pf_pipe1(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_pf_pipe2(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_pf_pipe3(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_pf_pipe4(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_pf_pipe5(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_pf_pipe6(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_pf_pipe7(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_ph_pipe0(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_ph_pipe1(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_ph_pipe2(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_ph_pipe3(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_ph_pipe4(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_ph_pipe5(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_ph_pipe6(),	 // Templated
		       .reg_rd_resv_pkt_cnt_lp_ph_pipe7(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fe_pipe0(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fe_pipe1(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fe_pipe2(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fe_pipe3(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fe_pipe4(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fe_pipe5(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fe_pipe6(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fe_pipe7(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fs_pipe0(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fs_pipe1(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fs_pipe2(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fs_pipe3(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fs_pipe4(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fs_pipe5(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fs_pipe6(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_fs_pipe7(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_le_pipe0(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_le_pipe1(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_le_pipe2(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_le_pipe3(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_le_pipe4(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_le_pipe5(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_le_pipe6(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_le_pipe7(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_ls_pipe0(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_ls_pipe1(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_ls_pipe2(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_ls_pipe3(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_ls_pipe4(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_ls_pipe5(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_ls_pipe6(),	 // Templated
		       .reg_rd_resv_pkt_cnt_sp_ls_pipe7(),	 // Templated
		       .reg_rd_send_pkt_cnt_lp_pf_aggr0(),	 // Templated
		       .reg_rd_send_pkt_cnt_lp_pf_aggr1(),	 // Templated
		       .reg_rd_send_pkt_cnt_lp_pf_aggr2(),	 // Templated
		       .reg_rd_send_pkt_cnt_lp_pf_aggr3(),	 // Templated
		       .reg_rd_send_pkt_cnt_lp_ph_aggr0(),	 // Templated
		       .reg_rd_send_pkt_cnt_lp_ph_aggr1(),	 // Templated
		       .reg_rd_send_pkt_cnt_lp_ph_aggr2(),	 // Templated
		       .reg_rd_send_pkt_cnt_lp_ph_aggr3(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_fe_aggr0(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_fe_aggr1(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_fe_aggr2(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_fe_aggr3(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_fs_aggr0(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_fs_aggr1(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_fs_aggr2(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_fs_aggr3(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_le_aggr0(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_le_aggr1(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_le_aggr2(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_le_aggr3(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_ls_aggr0(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_ls_aggr1(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_ls_aggr2(),	 // Templated
		       .reg_rd_send_pkt_cnt_sp_ls_aggr3(),	 // Templated
		       .reg_rd_vprbs_rx_check_app_route_lane0(), // Templated
		       .reg_rd_vprbs_rx_check_app_route_lane1(), // Templated
		       .reg_rd_vprbs_rx_check_app_route_lane2(), // Templated
		       .reg_rd_vprbs_rx_check_app_route_lane3(), // Templated
		       .reg_rd_vprbs_rx_check_app_route_lane4(), // Templated
		       .reg_rd_vprbs_rx_check_app_route_lane5(), // Templated
		       .reg_rd_vprbs_rx_check_app_route_lane6(), // Templated
		       .reg_rd_vprbs_rx_check_app_route_lane7(), // Templated
		       .reg_rd_vprbs_rx_err_app_route_lane0(),	 // Templated
		       .reg_rd_vprbs_rx_err_app_route_lane1(),	 // Templated
		       .reg_rd_vprbs_rx_err_app_route_lane2(),	 // Templated
		       .reg_rd_vprbs_rx_err_app_route_lane3(),	 // Templated
		       .reg_rd_vprbs_rx_err_app_route_lane4(),	 // Templated
		       .reg_rd_vprbs_rx_err_app_route_lane5(),	 // Templated
		       .reg_rd_vprbs_rx_err_app_route_lane6(),	 // Templated
		       .reg_rd_vprbs_rx_err_app_route_lane7(),	 // Templated
		       .reg_rd_vprbs_rx_fail_app_route_lane0(),	 // Templated
		       .reg_rd_vprbs_rx_fail_app_route_lane1(),	 // Templated
		       .reg_rd_vprbs_rx_fail_app_route_lane2(),	 // Templated
		       .reg_rd_vprbs_rx_fail_app_route_lane3(),	 // Templated
		       .reg_rd_vprbs_rx_fail_app_route_lane4(),	 // Templated
		       .reg_rd_vprbs_rx_fail_app_route_lane5(),	 // Templated
		       .reg_rd_vprbs_rx_fail_app_route_lane6(),	 // Templated
		       .reg_rd_vprbs_rx_fail_app_route_lane7(),	 // Templated
		       .video_data_afifo_ecc_fault0(video_data_afifo_ecc_fault0),
		       .video_data_afifo_ecc_fault1(video_data_afifo_ecc_fault1),
		       .video_data_afifo_ecc_fault2(video_data_afifo_ecc_fault2),
		       .video_data_afifo_ecc_fault3(video_data_afifo_ecc_fault3),
		       .video_data_afifo_ecc_fault4(video_data_afifo_ecc_fault4),
		       .video_data_afifo_ecc_fault5(video_data_afifo_ecc_fault5),
		       .video_data_afifo_ecc_fault6(video_data_afifo_ecc_fault6),
		       .video_data_afifo_ecc_fault7(video_data_afifo_ecc_fault7),
		       .video_data_fwft_fifo_ecc_fault0(video_data_fwft_fifo_ecc_fault0),
		       .video_data_fwft_fifo_ecc_fault1(video_data_fwft_fifo_ecc_fault1),
		       .video_data_fwft_fifo_ecc_fault2(video_data_fwft_fifo_ecc_fault2),
		       .video_data_fwft_fifo_ecc_fault3(video_data_fwft_fifo_ecc_fault3),
		       .video_data_fwft_fifo_ecc_fault4(video_data_fwft_fifo_ecc_fault4),
		       .video_data_fwft_fifo_ecc_fault5(video_data_fwft_fifo_ecc_fault5),
		       .video_data_fwft_fifo_ecc_fault6(video_data_fwft_fifo_ecc_fault6),
		       .video_data_fwft_fifo_ecc_fault7(video_data_fwft_fifo_ecc_fault7),
		       .to_clkgen_fifo_wrclk_sel0(),		 // Templated
		       .to_clkgen_fifo_wrclk_sel1(),		 // Templated
		       .to_clkgen_fifo_wrclk_sel2(),		 // Templated
		       .to_clkgen_fifo_wrclk_sel3(),		 // Templated
		       .to_clkgen_fifo_wrclk_sel4(),		 // Templated
		       .to_clkgen_fifo_wrclk_sel5(),		 // Templated
		       .to_clkgen_fifo_wrclk_sel6(),		 // Templated
		       .to_clkgen_fifo_wrclk_sel7(),		 // Templated
		       .to_clkgen_fifo_rdclk_sel0(),		 // Templated
		       .to_clkgen_fifo_rdclk_sel1(),		 // Templated
		       .to_clkgen_fifo_rdclk_sel2(),		 // Templated
		       .to_clkgen_fifo_rdclk_sel3(),		 // Templated
		       .to_clkgen_fifo_rdclk_sel4(),		 // Templated
		       .to_clkgen_fifo_rdclk_sel5(),		 // Templated
		       .to_clkgen_fifo_rdclk_sel6(),		 // Templated
		       .to_clkgen_fifo_rdclk_sel7(),		 // Templated
		       .reg_rd_video_lock0(reg_rd_video_lock0),
		       .reg_rd_video_lock1(reg_rd_video_lock1),
		       .reg_rd_video_lock2(reg_rd_video_lock2),
		       .reg_rd_video_lock3(reg_rd_video_lock3),
		       .reg_rd_video_lock4(reg_rd_video_lock4),
		       .reg_rd_video_lock5(reg_rd_video_lock5),
		       .reg_rd_video_lock6(reg_rd_video_lock6),
		       .reg_rd_video_lock7(reg_rd_video_lock7),
		       .reg_rd_video_loss0(reg_rd_video_loss0),
		       .reg_rd_video_loss1(reg_rd_video_loss1),
		       .reg_rd_video_loss2(reg_rd_video_loss2),
		       .reg_rd_video_loss3(reg_rd_video_loss3),
		       .reg_rd_video_loss4(reg_rd_video_loss4),
		       .reg_rd_video_loss5(reg_rd_video_loss5),
		       .reg_rd_video_loss6(reg_rd_video_loss6),
		       .reg_rd_video_loss7(reg_rd_video_loss7),
		       .video_loss0	(video_loss0),
		       .video_loss1	(video_loss1),
		       .video_loss2	(video_loss2),
		       .video_loss3	(video_loss3),
		       .video_loss4	(video_loss4),
		       .video_loss5	(video_loss5),
		       .video_loss6	(video_loss6),
		       .video_loss7	(video_loss7),
		       .reg_rd_fifo_rd_ctrl_cs0(),		 // Templated
		       .reg_rd_fifo_rd_ctrl_cs1(),		 // Templated
		       .reg_rd_fifo_rd_ctrl_cs2(),		 // Templated
		       .reg_rd_fifo_rd_ctrl_cs3(),		 // Templated
		       .reg_rd_fifo_rd_ctrl_cs4(),		 // Templated
		       .reg_rd_fifo_rd_ctrl_cs5(),		 // Templated
		       .reg_rd_fifo_rd_ctrl_cs6(),		 // Templated
		       .reg_rd_fifo_rd_ctrl_cs7(),		 // Templated
		       .reg_rd_fs_detect_pipe0(reg_rd_fs_detect_pipe0),
		       .reg_rd_fs_detect_pipe1(reg_rd_fs_detect_pipe1),
		       .reg_rd_fs_detect_pipe2(reg_rd_fs_detect_pipe2),
		       .reg_rd_fs_detect_pipe3(reg_rd_fs_detect_pipe3),
		       .reg_rd_fs_detect_pipe4(reg_rd_fs_detect_pipe4),
		       .reg_rd_fs_detect_pipe5(reg_rd_fs_detect_pipe5),
		       .reg_rd_fs_detect_pipe6(reg_rd_fs_detect_pipe6),
		       .reg_rd_fs_detect_pipe7(reg_rd_fs_detect_pipe7),
		       .reg_rd_fs_cnt_pipe0(),			 // Templated
		       .reg_rd_fs_cnt_pipe1(),			 // Templated
		       .reg_rd_fs_cnt_pipe2(),			 // Templated
		       .reg_rd_fs_cnt_pipe3(),			 // Templated
		       .reg_rd_fs_cnt_pipe4(),			 // Templated
		       .reg_rd_fs_cnt_pipe5(),			 // Templated
		       .reg_rd_fs_cnt_pipe6(),			 // Templated
		       .reg_rd_fs_cnt_pipe7(),			 // Templated
		       .reg_rd_cnt_line_end_rd_side0(),		 // Templated
		       .reg_rd_cnt_line_end_rd_side1(),		 // Templated
		       .reg_rd_cnt_line_end_rd_side2(),		 // Templated
		       .reg_rd_cnt_line_end_rd_side3(),		 // Templated
		       .reg_rd_cnt_line_end_rd_side4(),		 // Templated
		       .reg_rd_cnt_line_end_rd_side5(),		 // Templated
		       .reg_rd_cnt_line_end_rd_side6(),		 // Templated
		       .reg_rd_cnt_line_end_rd_side7(),		 // Templated
		       .reg_rd_sch0_cs	(),			 // Templated
		       .reg_rd_sch1_cs	(),			 // Templated
		       .reg_rd_sch2_cs	(),			 // Templated
		       .reg_rd_sch3_cs	(),			 // Templated
		       .reg_rd_sch2post_video_data_vld0(reg_rd_sch2post_video_data_vld0),
		       .reg_rd_sch2post_video_data_vld1(reg_rd_sch2post_video_data_vld1),
		       .reg_rd_sch2post_video_data_vld2(reg_rd_sch2post_video_data_vld2),
		       .reg_rd_sch2post_video_data_vld3(reg_rd_sch2post_video_data_vld3),
		       .reg_rd_pipe2sch_video_data_vld0(reg_rd_pipe2sch_video_data_vld0),
		       .reg_rd_pipe2sch_video_data_vld1(reg_rd_pipe2sch_video_data_vld1),
		       .reg_rd_pipe2sch_video_data_vld2(reg_rd_pipe2sch_video_data_vld2),
		       .reg_rd_pipe2sch_video_data_vld3(reg_rd_pipe2sch_video_data_vld3),
		       .reg_rd_pipe2sch_video_data_vld4(reg_rd_pipe2sch_video_data_vld4),
		       .reg_rd_pipe2sch_video_data_vld5(reg_rd_pipe2sch_video_data_vld5),
		       .reg_rd_pipe2sch_video_data_vld6(reg_rd_pipe2sch_video_data_vld6),
		       .reg_rd_pipe2sch_video_data_vld7(reg_rd_pipe2sch_video_data_vld7),
		       .reg_rd_pipe0_dispatched_cnt_ready_for_sch(reg_rd_pipe0_dispatched_cnt_ready_for_sch[31:0]),
		       .reg_rd_pipe1_dispatched_cnt_ready_for_sch(reg_rd_pipe1_dispatched_cnt_ready_for_sch[31:0]),
		       .reg_rd_pipe2_dispatched_cnt_ready_for_sch(reg_rd_pipe2_dispatched_cnt_ready_for_sch[31:0]),
		       .reg_rd_pipe3_dispatched_cnt_ready_for_sch(reg_rd_pipe3_dispatched_cnt_ready_for_sch[31:0]),
		       .reg_rd_pipe4_dispatched_cnt_ready_for_sch(reg_rd_pipe4_dispatched_cnt_ready_for_sch[31:0]),
		       .reg_rd_pipe5_dispatched_cnt_ready_for_sch(reg_rd_pipe5_dispatched_cnt_ready_for_sch[31:0]),
		       .reg_rd_pipe6_dispatched_cnt_ready_for_sch(reg_rd_pipe6_dispatched_cnt_ready_for_sch[31:0]),
		       .reg_rd_pipe7_dispatched_cnt_ready_for_sch(reg_rd_pipe7_dispatched_cnt_ready_for_sch[31:0]),
		       .video_data_afifo_mem_double_err0(video_data_afifo_mem_double_err0),
		       .video_data_afifo_mem_double_err1(video_data_afifo_mem_double_err1),
		       .video_data_afifo_mem_double_err2(video_data_afifo_mem_double_err2),
		       .video_data_afifo_mem_double_err3(video_data_afifo_mem_double_err3),
		       .video_data_afifo_mem_double_err4(video_data_afifo_mem_double_err4),
		       .video_data_afifo_mem_double_err5(video_data_afifo_mem_double_err5),
		       .video_data_afifo_mem_double_err6(video_data_afifo_mem_double_err6),
		       .video_data_afifo_mem_double_err7(video_data_afifo_mem_double_err7),
		       .video_data_afifo_mem_single_err0(video_data_afifo_mem_single_err0),
		       .video_data_afifo_mem_single_err1(video_data_afifo_mem_single_err1),
		       .video_data_afifo_mem_single_err2(video_data_afifo_mem_single_err2),
		       .video_data_afifo_mem_single_err3(video_data_afifo_mem_single_err3),
		       .video_data_afifo_mem_single_err4(video_data_afifo_mem_single_err4),
		       .video_data_afifo_mem_single_err5(video_data_afifo_mem_single_err5),
		       .video_data_afifo_mem_single_err6(video_data_afifo_mem_single_err6),
		       .video_data_afifo_mem_single_err7(video_data_afifo_mem_single_err7),
		       .video_data_afifo_ovf_int0(video_data_afifo_ovf_int0), // Templated
		       .video_data_afifo_ovf_int1(video_data_afifo_ovf_int1), // Templated
		       .video_data_afifo_ovf_int2(video_data_afifo_ovf_int2), // Templated
		       .video_data_afifo_ovf_int3(video_data_afifo_ovf_int3), // Templated
		       .video_data_afifo_ovf_int4(video_data_afifo_ovf_int4), // Templated
		       .video_data_afifo_ovf_int5(video_data_afifo_ovf_int5), // Templated
		       .video_data_afifo_ovf_int6(video_data_afifo_ovf_int6), // Templated
		       .video_data_afifo_ovf_int7(video_data_afifo_ovf_int7), // Templated
		       .video_data_fwft_fifo_mem_double_err0(video_data_fwft_fifo_mem_double_err0),
		       .video_data_fwft_fifo_mem_double_err1(video_data_fwft_fifo_mem_double_err1),
		       .video_data_fwft_fifo_mem_double_err2(video_data_fwft_fifo_mem_double_err2),
		       .video_data_fwft_fifo_mem_double_err3(video_data_fwft_fifo_mem_double_err3),
		       .video_data_fwft_fifo_mem_double_err4(video_data_fwft_fifo_mem_double_err4),
		       .video_data_fwft_fifo_mem_double_err5(video_data_fwft_fifo_mem_double_err5),
		       .video_data_fwft_fifo_mem_double_err6(video_data_fwft_fifo_mem_double_err6),
		       .video_data_fwft_fifo_mem_double_err7(video_data_fwft_fifo_mem_double_err7),
		       .video_data_fwft_fifo_mem_single_err0(video_data_fwft_fifo_mem_single_err0),
		       .video_data_fwft_fifo_mem_single_err1(video_data_fwft_fifo_mem_single_err1),
		       .video_data_fwft_fifo_mem_single_err2(video_data_fwft_fifo_mem_single_err2),
		       .video_data_fwft_fifo_mem_single_err3(video_data_fwft_fifo_mem_single_err3),
		       .video_data_fwft_fifo_mem_single_err4(video_data_fwft_fifo_mem_single_err4),
		       .video_data_fwft_fifo_mem_single_err5(video_data_fwft_fifo_mem_single_err5),
		       .video_data_fwft_fifo_mem_single_err6(video_data_fwft_fifo_mem_single_err6),
		       .video_data_fwft_fifo_mem_single_err7(video_data_fwft_fifo_mem_single_err7),
		       .video_data_fwft_fifo_ovf_int0(video_data_fwft_fifo_ovf_int0),
		       .video_data_fwft_fifo_ovf_int1(video_data_fwft_fifo_ovf_int1),
		       .video_data_fwft_fifo_ovf_int2(video_data_fwft_fifo_ovf_int2),
		       .video_data_fwft_fifo_ovf_int3(video_data_fwft_fifo_ovf_int3),
		       .video_data_fwft_fifo_ovf_int4(video_data_fwft_fifo_ovf_int4),
		       .video_data_fwft_fifo_ovf_int5(video_data_fwft_fifo_ovf_int5),
		       .video_data_fwft_fifo_ovf_int6(video_data_fwft_fifo_ovf_int6),
		       .video_data_fwft_fifo_ovf_int7(video_data_fwft_fifo_ovf_int7),
		       .lcrc_err0	(lcrc_err0),
		       .lcrc_err1	(lcrc_err1),
		       .lcrc_err2	(lcrc_err2),
		       .lcrc_err3	(lcrc_err3),
		       .lcrc_err4	(lcrc_err4),
		       .lcrc_err5	(lcrc_err5),
		       .lcrc_err6	(lcrc_err6),
		       .lcrc_err7	(lcrc_err7),
		       .vprbs_rx_fail_app_route_int0(),		 // Templated
		       .vprbs_rx_fail_app_route_int1(),		 // Templated
		       .vprbs_rx_fail_app_route_int2(),		 // Templated
		       .vprbs_rx_fail_app_route_int3(),		 // Templated
		       .vprbs_rx_fail_app_route_int4(),		 // Templated
		       .vprbs_rx_fail_app_route_int5(),		 // Templated
		       .vprbs_rx_fail_app_route_int6(),		 // Templated
		       .vprbs_rx_fail_app_route_int7(),		 // Templated
		       .sch_data_type_align_fail_int0(sch_data_type_align_fail_int0),
		       .sch_data_type_align_fail_int1(sch_data_type_align_fail_int1),
		       .sch_data_type_align_fail_int2(sch_data_type_align_fail_int2),
		       .sch_data_type_align_fail_int3(sch_data_type_align_fail_int3),
		       // Inputs
		       .aggre_clk0	(aggre_clk0),
		       .aggre_clk1	(aggre_clk1),
		       .aggre_clk2	(aggre_clk2),
		       .aggre_clk3	(aggre_clk3),
		       .aggre_clk_rst_n0(aggre_clk_rst_n0),
		       .aggre_clk_rst_n1(aggre_clk_rst_n1),
		       .aggre_clk_rst_n2(aggre_clk_rst_n2),
		       .aggre_clk_rst_n3(aggre_clk_rst_n3),
		       .clk_1M		(clk_1M),
		       .clk_1M_rst_n	(clk_1M_rst_n),
		       .fifo_rdclk0	(fifo_rdclk0),
		       .fifo_rdclk1	(fifo_rdclk1),
		       .fifo_rdclk2	(fifo_rdclk2),
		       .fifo_rdclk3	(fifo_rdclk3),
		       .fifo_rdclk4	(fifo_rdclk4),
		       .fifo_rdclk5	(fifo_rdclk5),
		       .fifo_rdclk6	(fifo_rdclk6),
		       .fifo_rdclk7	(fifo_rdclk7),
		       .fifo_rdclk_rst_n0(fifo_rdclk_rst_n0),
		       .fifo_rdclk_rst_n1(fifo_rdclk_rst_n1),
		       .fifo_rdclk_rst_n2(fifo_rdclk_rst_n2),
		       .fifo_rdclk_rst_n3(fifo_rdclk_rst_n3),
		       .fifo_rdclk_rst_n4(fifo_rdclk_rst_n4),
		       .fifo_rdclk_rst_n5(fifo_rdclk_rst_n5),
		       .fifo_rdclk_rst_n6(fifo_rdclk_rst_n6),
		       .fifo_rdclk_rst_n7(fifo_rdclk_rst_n7),
		       .fifo_wrclk0	(fifo_wrclk0),
		       .fifo_wrclk1	(fifo_wrclk1),
		       .fifo_wrclk2	(fifo_wrclk2),
		       .fifo_wrclk3	(fifo_wrclk3),
		       .fifo_wrclk4	(fifo_wrclk4),
		       .fifo_wrclk5	(fifo_wrclk5),
		       .fifo_wrclk6	(fifo_wrclk6),
		       .fifo_wrclk7	(fifo_wrclk7),
		       .fifo_wrclk_rst_n0(fifo_wrclk_rst_n0),
		       .fifo_wrclk_rst_n1(fifo_wrclk_rst_n1),
		       .fifo_wrclk_rst_n2(fifo_wrclk_rst_n2),
		       .fifo_wrclk_rst_n3(fifo_wrclk_rst_n3),
		       .fifo_wrclk_rst_n4(fifo_wrclk_rst_n4),
		       .fifo_wrclk_rst_n5(fifo_wrclk_rst_n5),
		       .fifo_wrclk_rst_n6(fifo_wrclk_rst_n6),
		       .fifo_wrclk_rst_n7(fifo_wrclk_rst_n7),
		       .gpio2app_sch0_frame_sync_lock(gpio2app_sch0_frame_sync_lock),
		       .gpio2app_sch1_frame_sync_lock(gpio2app_sch1_frame_sync_lock),
		       .gpio2app_sch2_frame_sync_lock(gpio2app_sch2_frame_sync_lock),
		       .gpio2app_sch3_frame_sync_lock(gpio2app_sch3_frame_sync_lock),
		       .mep0_byte_en	(idi_byte_en_lane0[2:0]), // Templated
		       .mep0_csi_data	(idi_data_lane0[63:0]),	 // Templated
		       .mep0_data_en	(idi_data_en_lane0),	 // Templated
		       .mep0_data_type	(idi_dt_lane0[5:0]),	 // Templated
		       .mep0_header_en	(idi_header_en_lane0),	 // Templated
		       .mep0_tunnel_mode_en(1'd0),		 // Templated
		       .mep0_word_count	(idi_word_count_lane0[15:0]), // Templated
		       .mep1_byte_en	(idi_byte_en_lane1[2:0]), // Templated
		       .mep1_csi_data	(idi_data_lane1[63:0]),	 // Templated
		       .mep1_data_en	(idi_data_en_lane1),	 // Templated
		       .mep1_data_type	(idi_dt_lane1[5:0]),	 // Templated
		       .mep1_header_en	(idi_header_en_lane1),	 // Templated
		       .mep1_tunnel_mode_en(1'd0),		 // Templated
		       .mep1_word_count	(idi_word_count_lane1[15:0]), // Templated
		       .mep2_byte_en	(idi_byte_en_lane2[2:0]), // Templated
		       .mep2_csi_data	(idi_data_lane2[63:0]),	 // Templated
		       .mep2_data_en	(idi_data_en_lane2),	 // Templated
		       .mep2_data_type	(idi_dt_lane2[5:0]),	 // Templated
		       .mep2_header_en	(idi_header_en_lane2),	 // Templated
		       .mep2_tunnel_mode_en(1'd0),		 // Templated
		       .mep2_word_count	(idi_word_count_lane2[15:0]), // Templated
		       .mep3_byte_en	(idi_byte_en_lane3[2:0]), // Templated
		       .mep3_csi_data	(idi_data_lane3[63:0]),	 // Templated
		       .mep3_data_en	(idi_data_en_lane3),	 // Templated
		       .mep3_data_type	(idi_dt_lane3[5:0]),	 // Templated
		       .mep3_header_en	(idi_header_en_lane3),	 // Templated
		       .mep3_tunnel_mode_en(1'd0),		 // Templated
		       .mep3_word_count	(idi_word_count_lane3[15:0]), // Templated
		       .reg_all_pipe_wr_mode_strobe(reg_all_pipe_wr_mode_strobe),
		       .reg_app_aggr0_vc_bit_override_en(reg_app_aggr0_vc_bit_override_en[2:0]),
		       .reg_app_aggr0_vc_bit_override_value(reg_app_aggr0_vc_bit_override_value[2:0]),
		       .reg_app_aggr1_vc_bit_override_en(reg_app_aggr1_vc_bit_override_en[2:0]),
		       .reg_app_aggr1_vc_bit_override_value(reg_app_aggr1_vc_bit_override_value[2:0]),
		       .reg_app_aggr2_vc_bit_override_en(reg_app_aggr2_vc_bit_override_en[2:0]),
		       .reg_app_aggr2_vc_bit_override_value(reg_app_aggr2_vc_bit_override_value[2:0]),
		       .reg_app_aggr3_vc_bit_override_en(reg_app_aggr3_vc_bit_override_en[2:0]),
		       .reg_app_aggr3_vc_bit_override_value(reg_app_aggr3_vc_bit_override_value[2:0]),
		       .reg_app_aggr_idi_crc_chk_en(reg_app_aggr_idi_crc_chk_en[3:0]),
		       .reg_app_ecc_addr_protect_en(1'd1),	 // Templated
		       .reg_app_ecc_bypass(1'd0),		 // Templated
		       .reg_app_ecc_fault_detc_en(1'd1),	 // Templated
		       .reg_app_pkt_crc_gen_dis(reg_app_pkt_crc_gen_dis),
		       .reg_app_sch0_frame_sync_lock(reg_app_sch0_frame_sync_lock),
		       .reg_app_sch0_frame_sync_lock_force(reg_app_sch0_frame_sync_lock_force),
		       .reg_app_sch1_frame_sync_lock(reg_app_sch1_frame_sync_lock),
		       .reg_app_sch1_frame_sync_lock_force(reg_app_sch1_frame_sync_lock_force),
		       .reg_app_sch2_frame_sync_lock(reg_app_sch2_frame_sync_lock),
		       .reg_app_sch2_frame_sync_lock_force(reg_app_sch2_frame_sync_lock_force),
		       .reg_app_sch3_frame_sync_lock(reg_app_sch3_frame_sync_lock),
		       .reg_app_sch3_frame_sync_lock_force(reg_app_sch3_frame_sync_lock_force),
		       .reg_app_wr_idi_data_continue(reg_app_wr_idi_data_continue),
		       .reg_clear_app_full_cnt_async_fifo_pipe0(reg_clear_app_full_cnt_async_fifo_pipe0),
		       .reg_clear_app_full_cnt_async_fifo_pipe1(reg_clear_app_full_cnt_async_fifo_pipe1),
		       .reg_clear_app_full_cnt_async_fifo_pipe2(reg_clear_app_full_cnt_async_fifo_pipe2),
		       .reg_clear_app_full_cnt_async_fifo_pipe3(reg_clear_app_full_cnt_async_fifo_pipe3),
		       .reg_clear_app_full_cnt_async_fifo_pipe4(reg_clear_app_full_cnt_async_fifo_pipe4),
		       .reg_clear_app_full_cnt_async_fifo_pipe5(reg_clear_app_full_cnt_async_fifo_pipe5),
		       .reg_clear_app_full_cnt_async_fifo_pipe6(reg_clear_app_full_cnt_async_fifo_pipe6),
		       .reg_clear_app_full_cnt_async_fifo_pipe7(reg_clear_app_full_cnt_async_fifo_pipe7),
		       .reg_clear_app_full_cnt_sync_fifo_pipe0(reg_clear_app_full_cnt_sync_fifo_pipe0),
		       .reg_clear_app_full_cnt_sync_fifo_pipe1(reg_clear_app_full_cnt_sync_fifo_pipe1),
		       .reg_clear_app_full_cnt_sync_fifo_pipe2(reg_clear_app_full_cnt_sync_fifo_pipe2),
		       .reg_clear_app_full_cnt_sync_fifo_pipe3(reg_clear_app_full_cnt_sync_fifo_pipe3),
		       .reg_clear_app_full_cnt_sync_fifo_pipe4(reg_clear_app_full_cnt_sync_fifo_pipe4),
		       .reg_clear_app_full_cnt_sync_fifo_pipe5(reg_clear_app_full_cnt_sync_fifo_pipe5),
		       .reg_clear_app_full_cnt_sync_fifo_pipe6(reg_clear_app_full_cnt_sync_fifo_pipe6),
		       .reg_clear_app_full_cnt_sync_fifo_pipe7(reg_clear_app_full_cnt_sync_fifo_pipe7),
		       .reg_clear_resv_pkt_cnt_lp_pf_pipe0(reg_clear_resv_pkt_cnt_lp_pf), // Templated
		       .reg_clear_resv_pkt_cnt_lp_pf_pipe1(reg_clear_resv_pkt_cnt_lp_pf), // Templated
		       .reg_clear_resv_pkt_cnt_lp_pf_pipe2(reg_clear_resv_pkt_cnt_lp_pf), // Templated
		       .reg_clear_resv_pkt_cnt_lp_pf_pipe3(reg_clear_resv_pkt_cnt_lp_pf), // Templated
		       .reg_clear_resv_pkt_cnt_lp_pf_pipe4(reg_clear_resv_pkt_cnt_lp_pf), // Templated
		       .reg_clear_resv_pkt_cnt_lp_pf_pipe5(reg_clear_resv_pkt_cnt_lp_pf), // Templated
		       .reg_clear_resv_pkt_cnt_lp_pf_pipe6(reg_clear_resv_pkt_cnt_lp_pf), // Templated
		       .reg_clear_resv_pkt_cnt_lp_pf_pipe7(reg_clear_resv_pkt_cnt_lp_pf), // Templated
		       .reg_clear_resv_pkt_cnt_lp_ph_pipe0(reg_clear_resv_pkt_cnt_lp_ph), // Templated
		       .reg_clear_resv_pkt_cnt_lp_ph_pipe1(reg_clear_resv_pkt_cnt_lp_ph), // Templated
		       .reg_clear_resv_pkt_cnt_lp_ph_pipe2(reg_clear_resv_pkt_cnt_lp_ph), // Templated
		       .reg_clear_resv_pkt_cnt_lp_ph_pipe3(reg_clear_resv_pkt_cnt_lp_ph), // Templated
		       .reg_clear_resv_pkt_cnt_lp_ph_pipe4(reg_clear_resv_pkt_cnt_lp_ph), // Templated
		       .reg_clear_resv_pkt_cnt_lp_ph_pipe5(reg_clear_resv_pkt_cnt_lp_ph), // Templated
		       .reg_clear_resv_pkt_cnt_lp_ph_pipe6(reg_clear_resv_pkt_cnt_lp_ph), // Templated
		       .reg_clear_resv_pkt_cnt_lp_ph_pipe7(reg_clear_resv_pkt_cnt_lp_ph), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fe_pipe0(reg_clear_resv_pkt_cnt_sp_fe), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fe_pipe1(reg_clear_resv_pkt_cnt_sp_fe), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fe_pipe2(reg_clear_resv_pkt_cnt_sp_fe), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fe_pipe3(reg_clear_resv_pkt_cnt_sp_fe), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fe_pipe4(reg_clear_resv_pkt_cnt_sp_fe), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fe_pipe5(reg_clear_resv_pkt_cnt_sp_fe), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fe_pipe6(reg_clear_resv_pkt_cnt_sp_fe), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fe_pipe7(reg_clear_resv_pkt_cnt_sp_fe), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fs_pipe0(reg_clear_resv_pkt_cnt_sp_fs), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fs_pipe1(reg_clear_resv_pkt_cnt_sp_fs), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fs_pipe2(reg_clear_resv_pkt_cnt_sp_fs), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fs_pipe3(reg_clear_resv_pkt_cnt_sp_fs), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fs_pipe4(reg_clear_resv_pkt_cnt_sp_fs), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fs_pipe5(reg_clear_resv_pkt_cnt_sp_fs), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fs_pipe6(reg_clear_resv_pkt_cnt_sp_fs), // Templated
		       .reg_clear_resv_pkt_cnt_sp_fs_pipe7(reg_clear_resv_pkt_cnt_sp_fs), // Templated
		       .reg_clear_resv_pkt_cnt_sp_le_pipe0(reg_clear_resv_pkt_cnt_sp_le), // Templated
		       .reg_clear_resv_pkt_cnt_sp_le_pipe1(reg_clear_resv_pkt_cnt_sp_le), // Templated
		       .reg_clear_resv_pkt_cnt_sp_le_pipe2(reg_clear_resv_pkt_cnt_sp_le), // Templated
		       .reg_clear_resv_pkt_cnt_sp_le_pipe3(reg_clear_resv_pkt_cnt_sp_le), // Templated
		       .reg_clear_resv_pkt_cnt_sp_le_pipe4(reg_clear_resv_pkt_cnt_sp_le), // Templated
		       .reg_clear_resv_pkt_cnt_sp_le_pipe5(reg_clear_resv_pkt_cnt_sp_le), // Templated
		       .reg_clear_resv_pkt_cnt_sp_le_pipe6(reg_clear_resv_pkt_cnt_sp_le), // Templated
		       .reg_clear_resv_pkt_cnt_sp_le_pipe7(reg_clear_resv_pkt_cnt_sp_le), // Templated
		       .reg_clear_resv_pkt_cnt_sp_ls_pipe0(reg_clear_resv_pkt_cnt_sp_ls), // Templated
		       .reg_clear_resv_pkt_cnt_sp_ls_pipe1(reg_clear_resv_pkt_cnt_sp_ls), // Templated
		       .reg_clear_resv_pkt_cnt_sp_ls_pipe2(reg_clear_resv_pkt_cnt_sp_ls), // Templated
		       .reg_clear_resv_pkt_cnt_sp_ls_pipe3(reg_clear_resv_pkt_cnt_sp_ls), // Templated
		       .reg_clear_resv_pkt_cnt_sp_ls_pipe4(reg_clear_resv_pkt_cnt_sp_ls), // Templated
		       .reg_clear_resv_pkt_cnt_sp_ls_pipe5(reg_clear_resv_pkt_cnt_sp_ls), // Templated
		       .reg_clear_resv_pkt_cnt_sp_ls_pipe6(reg_clear_resv_pkt_cnt_sp_ls), // Templated
		       .reg_clear_resv_pkt_cnt_sp_ls_pipe7(reg_clear_resv_pkt_cnt_sp_ls), // Templated
		       .reg_clear_send_pkt_cnt_lp_pf_aggr0(reg_clear_send_pkt_cnt_lp_pf), // Templated
		       .reg_clear_send_pkt_cnt_lp_pf_aggr1(reg_clear_send_pkt_cnt_lp_pf), // Templated
		       .reg_clear_send_pkt_cnt_lp_pf_aggr2(reg_clear_send_pkt_cnt_lp_pf), // Templated
		       .reg_clear_send_pkt_cnt_lp_pf_aggr3(reg_clear_send_pkt_cnt_lp_pf), // Templated
		       .reg_clear_send_pkt_cnt_lp_ph_aggr0(reg_clear_send_pkt_cnt_lp_ph), // Templated
		       .reg_clear_send_pkt_cnt_lp_ph_aggr1(reg_clear_send_pkt_cnt_lp_ph), // Templated
		       .reg_clear_send_pkt_cnt_lp_ph_aggr2(reg_clear_send_pkt_cnt_lp_ph), // Templated
		       .reg_clear_send_pkt_cnt_lp_ph_aggr3(reg_clear_send_pkt_cnt_lp_ph), // Templated
		       .reg_clear_send_pkt_cnt_sp_fe_aggr0(reg_clear_send_pkt_cnt_sp_fe), // Templated
		       .reg_clear_send_pkt_cnt_sp_fe_aggr1(reg_clear_send_pkt_cnt_sp_fe), // Templated
		       .reg_clear_send_pkt_cnt_sp_fe_aggr2(reg_clear_send_pkt_cnt_sp_fe), // Templated
		       .reg_clear_send_pkt_cnt_sp_fe_aggr3(reg_clear_send_pkt_cnt_sp_fe), // Templated
		       .reg_clear_send_pkt_cnt_sp_fs_aggr0(reg_clear_send_pkt_cnt_sp_fs), // Templated
		       .reg_clear_send_pkt_cnt_sp_fs_aggr1(reg_clear_send_pkt_cnt_sp_fs), // Templated
		       .reg_clear_send_pkt_cnt_sp_fs_aggr2(reg_clear_send_pkt_cnt_sp_fs), // Templated
		       .reg_clear_send_pkt_cnt_sp_fs_aggr3(reg_clear_send_pkt_cnt_sp_fs), // Templated
		       .reg_clear_send_pkt_cnt_sp_le_aggr0(reg_clear_send_pkt_cnt_sp_le), // Templated
		       .reg_clear_send_pkt_cnt_sp_le_aggr1(reg_clear_send_pkt_cnt_sp_le), // Templated
		       .reg_clear_send_pkt_cnt_sp_le_aggr2(reg_clear_send_pkt_cnt_sp_le), // Templated
		       .reg_clear_send_pkt_cnt_sp_le_aggr3(reg_clear_send_pkt_cnt_sp_le), // Templated
		       .reg_clear_send_pkt_cnt_sp_ls_aggr0(reg_clear_send_pkt_cnt_sp_ls), // Templated
		       .reg_clear_send_pkt_cnt_sp_ls_aggr1(reg_clear_send_pkt_cnt_sp_ls), // Templated
		       .reg_clear_send_pkt_cnt_sp_ls_aggr2(reg_clear_send_pkt_cnt_sp_ls), // Templated
		       .reg_clear_send_pkt_cnt_sp_ls_aggr3(reg_clear_send_pkt_cnt_sp_ls), // Templated
		       .reg_dbg_pkt_num_nonzero_and_fifo_empty_threshold(16'd200), // Templated
		       .reg_dbg_pkt_num_nonzero_threshold(16'd200), // Templated
		       .reg_delete_lp_depend_on_wc_mux(reg_delete_lp_depend_on_wc_mux),
		       .reg_dft_sync_tpram_config(10'd0),	 // Templated
		       .reg_dft_tpram_config(9'd0),		 // Templated
		       .reg_drop_mapping_fault_pkt(reg_drop_mapping_fault_pkt[7:0]),
		       .reg_last_byte_header_down_mux(reg_last_byte_header_down_mux),
		       .reg_mem_dt1_selz_mep0(reg_mem_dt1_selz[6:0]), // Templated
		       .reg_mem_dt1_selz_mep1(reg_mem_dt1_selz[6:0]), // Templated
		       .reg_mem_dt1_selz_mep2(reg_mem_dt1_selz[6:0]), // Templated
		       .reg_mem_dt1_selz_mep3(reg_mem_dt1_selz[6:0]), // Templated
		       .reg_mem_dt2_selz_mep0(reg_mem_dt2_selz[6:0]), // Templated
		       .reg_mem_dt2_selz_mep1(reg_mem_dt2_selz[6:0]), // Templated
		       .reg_mem_dt2_selz_mep2(reg_mem_dt2_selz[6:0]), // Templated
		       .reg_mem_dt2_selz_mep3(reg_mem_dt2_selz[6:0]), // Templated
		       .reg_mem_dt3_selz_en_mep0(reg_mem_dt3_selz_en), // Templated
		       .reg_mem_dt3_selz_en_mep1(reg_mem_dt3_selz_en), // Templated
		       .reg_mem_dt3_selz_en_mep2(reg_mem_dt3_selz_en), // Templated
		       .reg_mem_dt3_selz_en_mep3(reg_mem_dt3_selz_en), // Templated
		       .reg_mem_dt3_selz_mep0(reg_mem_dt3_selz[7:0]), // Templated
		       .reg_mem_dt3_selz_mep1(reg_mem_dt3_selz[7:0]), // Templated
		       .reg_mem_dt3_selz_mep2(reg_mem_dt3_selz[7:0]), // Templated
		       .reg_mem_dt3_selz_mep3(reg_mem_dt3_selz[7:0]), // Templated
		       .reg_mem_dt4_selz_en_mep0(reg_mem_dt4_selz_en), // Templated
		       .reg_mem_dt4_selz_en_mep1(reg_mem_dt4_selz_en), // Templated
		       .reg_mem_dt4_selz_en_mep2(reg_mem_dt4_selz_en), // Templated
		       .reg_mem_dt4_selz_en_mep3(reg_mem_dt4_selz_en), // Templated
		       .reg_mem_dt4_selz_mep0(reg_mem_dt4_selz[7:0]), // Templated
		       .reg_mem_dt4_selz_mep1(reg_mem_dt4_selz[7:0]), // Templated
		       .reg_mem_dt4_selz_mep2(reg_mem_dt4_selz[7:0]), // Templated
		       .reg_mem_dt4_selz_mep3(reg_mem_dt4_selz[7:0]), // Templated
		       .reg_mem_dt7_selz_mep0(reg_mem_dt7_selz[6:0]), // Templated
		       .reg_mem_dt7_selz_mep1(reg_mem_dt7_selz[6:0]), // Templated
		       .reg_mem_dt7_selz_mep2(reg_mem_dt7_selz[6:0]), // Templated
		       .reg_mem_dt7_selz_mep3(reg_mem_dt7_selz[6:0]), // Templated
		       .reg_mem_dt8_selz_mep0(reg_mem_dt8_selz[6:0]), // Templated
		       .reg_mem_dt8_selz_mep1(reg_mem_dt8_selz[6:0]), // Templated
		       .reg_mem_dt8_selz_mep2(reg_mem_dt8_selz[6:0]), // Templated
		       .reg_mem_dt8_selz_mep3(reg_mem_dt8_selz[6:0]), // Templated
		       .reg_mep0_tdi_en	(1'd0),			 // Templated
		       .reg_mep0_tdi_en_force(1'd0),		 // Templated
		       .reg_mep1_tdi_en	(1'd0),			 // Templated
		       .reg_mep1_tdi_en_force(1'd0),		 // Templated
		       .reg_mep2_tdi_en	(1'd0),			 // Templated
		       .reg_mep2_tdi_en_force(1'd0),		 // Templated
		       .reg_mep3_tdi_en	(1'd0),			 // Templated
		       .reg_mep3_tdi_en_force(1'd0),		 // Templated
		       .reg_pipe0_drop_ls_le_pkt(reg_pipe0_drop_ls_le_pkt),
		       .reg_pipe0_map0_aggr_id(reg_pipe0_map0_aggr_id), // Templated
		       .reg_pipe0_map0_dt_dest(reg_pipe0_map0_dt_dest ), // Templated
		       .reg_pipe0_map0_dt_source(reg_pipe0_map0_dt_source ), // Templated
		       .reg_pipe0_map0_vc_dest(reg_pipe0_map0_vc_dest ), // Templated
		       .reg_pipe0_map0_vc_source(reg_pipe0_map0_vc_source ), // Templated
		       .reg_pipe0_map10_aggr_id(reg_pipe0_map10_aggr_id), // Templated
		       .reg_pipe0_map10_dt_dest(reg_pipe0_map10_dt_dest), // Templated
		       .reg_pipe0_map10_dt_source(reg_pipe0_map10_dt_source), // Templated
		       .reg_pipe0_map10_vc_dest(reg_pipe0_map10_vc_dest), // Templated
		       .reg_pipe0_map10_vc_source(reg_pipe0_map10_vc_source), // Templated
		       .reg_pipe0_map11_aggr_id(reg_pipe0_map11_aggr_id), // Templated
		       .reg_pipe0_map11_dt_dest(reg_pipe0_map11_dt_dest), // Templated
		       .reg_pipe0_map11_dt_source(reg_pipe0_map11_dt_source), // Templated
		       .reg_pipe0_map11_vc_dest(reg_pipe0_map11_vc_dest), // Templated
		       .reg_pipe0_map11_vc_source(reg_pipe0_map11_vc_source), // Templated
		       .reg_pipe0_map12_aggr_id(reg_pipe0_map12_aggr_id), // Templated
		       .reg_pipe0_map12_dt_dest(reg_pipe0_map12_dt_dest), // Templated
		       .reg_pipe0_map12_dt_source(reg_pipe0_map12_dt_source), // Templated
		       .reg_pipe0_map12_vc_dest(reg_pipe0_map12_vc_dest), // Templated
		       .reg_pipe0_map12_vc_source(reg_pipe0_map12_vc_source), // Templated
		       .reg_pipe0_map13_aggr_id(reg_pipe0_map13_aggr_id), // Templated
		       .reg_pipe0_map13_dt_dest(reg_pipe0_map13_dt_dest), // Templated
		       .reg_pipe0_map13_dt_source(reg_pipe0_map13_dt_source), // Templated
		       .reg_pipe0_map13_vc_dest(reg_pipe0_map13_vc_dest), // Templated
		       .reg_pipe0_map13_vc_source(reg_pipe0_map13_vc_source), // Templated
		       .reg_pipe0_map14_aggr_id(reg_pipe0_map14_aggr_id), // Templated
		       .reg_pipe0_map14_dt_dest(reg_pipe0_map14_dt_dest), // Templated
		       .reg_pipe0_map14_dt_source(reg_pipe0_map14_dt_source), // Templated
		       .reg_pipe0_map14_vc_dest(reg_pipe0_map14_vc_dest), // Templated
		       .reg_pipe0_map14_vc_source(reg_pipe0_map14_vc_source), // Templated
		       .reg_pipe0_map15_aggr_id(reg_pipe0_map15_aggr_id), // Templated
		       .reg_pipe0_map15_dt_dest(reg_pipe0_map15_dt_dest), // Templated
		       .reg_pipe0_map15_dt_source(reg_pipe0_map15_dt_source), // Templated
		       .reg_pipe0_map15_vc_dest(reg_pipe0_map15_vc_dest), // Templated
		       .reg_pipe0_map15_vc_source(reg_pipe0_map15_vc_source), // Templated
		       .reg_pipe0_map1_aggr_id(reg_pipe0_map1_aggr_id), // Templated
		       .reg_pipe0_map1_dt_dest(reg_pipe0_map1_dt_dest ), // Templated
		       .reg_pipe0_map1_dt_source(reg_pipe0_map1_dt_source ), // Templated
		       .reg_pipe0_map1_vc_dest(reg_pipe0_map1_vc_dest ), // Templated
		       .reg_pipe0_map1_vc_source(reg_pipe0_map1_vc_source ), // Templated
		       .reg_pipe0_map2_aggr_id(reg_pipe0_map2_aggr_id), // Templated
		       .reg_pipe0_map2_dt_dest(reg_pipe0_map2_dt_dest ), // Templated
		       .reg_pipe0_map2_dt_source(reg_pipe0_map2_dt_source ), // Templated
		       .reg_pipe0_map2_vc_dest(reg_pipe0_map2_vc_dest ), // Templated
		       .reg_pipe0_map2_vc_source(reg_pipe0_map2_vc_source ), // Templated
		       .reg_pipe0_map3_aggr_id(reg_pipe0_map3_aggr_id), // Templated
		       .reg_pipe0_map3_dt_dest(reg_pipe0_map3_dt_dest ), // Templated
		       .reg_pipe0_map3_dt_source(reg_pipe0_map3_dt_source ), // Templated
		       .reg_pipe0_map3_vc_dest(reg_pipe0_map3_vc_dest ), // Templated
		       .reg_pipe0_map3_vc_source(reg_pipe0_map3_vc_source ), // Templated
		       .reg_pipe0_map4_aggr_id(reg_pipe0_map4_aggr_id), // Templated
		       .reg_pipe0_map4_dt_dest(reg_pipe0_map4_dt_dest ), // Templated
		       .reg_pipe0_map4_dt_source(reg_pipe0_map4_dt_source ), // Templated
		       .reg_pipe0_map4_vc_dest(reg_pipe0_map4_vc_dest ), // Templated
		       .reg_pipe0_map4_vc_source(reg_pipe0_map4_vc_source ), // Templated
		       .reg_pipe0_map5_aggr_id(reg_pipe0_map5_aggr_id), // Templated
		       .reg_pipe0_map5_dt_dest(reg_pipe0_map5_dt_dest ), // Templated
		       .reg_pipe0_map5_dt_source(reg_pipe0_map5_dt_source ), // Templated
		       .reg_pipe0_map5_vc_dest(reg_pipe0_map5_vc_dest ), // Templated
		       .reg_pipe0_map5_vc_source(reg_pipe0_map5_vc_source ), // Templated
		       .reg_pipe0_map6_aggr_id(reg_pipe0_map6_aggr_id), // Templated
		       .reg_pipe0_map6_dt_dest(reg_pipe0_map6_dt_dest ), // Templated
		       .reg_pipe0_map6_dt_source(reg_pipe0_map6_dt_source ), // Templated
		       .reg_pipe0_map6_vc_dest(reg_pipe0_map6_vc_dest ), // Templated
		       .reg_pipe0_map6_vc_source(reg_pipe0_map6_vc_source ), // Templated
		       .reg_pipe0_map7_aggr_id(reg_pipe0_map7_aggr_id), // Templated
		       .reg_pipe0_map7_dt_dest(reg_pipe0_map7_dt_dest ), // Templated
		       .reg_pipe0_map7_dt_source(reg_pipe0_map7_dt_source ), // Templated
		       .reg_pipe0_map7_vc_dest(reg_pipe0_map7_vc_dest ), // Templated
		       .reg_pipe0_map7_vc_source(reg_pipe0_map7_vc_source ), // Templated
		       .reg_pipe0_map8_aggr_id(reg_pipe0_map8_aggr_id), // Templated
		       .reg_pipe0_map8_dt_dest(reg_pipe0_map8_dt_dest ), // Templated
		       .reg_pipe0_map8_dt_source(reg_pipe0_map8_dt_source ), // Templated
		       .reg_pipe0_map8_vc_dest(reg_pipe0_map8_vc_dest ), // Templated
		       .reg_pipe0_map8_vc_source(reg_pipe0_map8_vc_source ), // Templated
		       .reg_pipe0_map9_aggr_id(reg_pipe0_map9_aggr_id), // Templated
		       .reg_pipe0_map9_dt_dest(reg_pipe0_map9_dt_dest ), // Templated
		       .reg_pipe0_map9_dt_source(reg_pipe0_map9_dt_source ), // Templated
		       .reg_pipe0_map9_vc_dest(reg_pipe0_map9_vc_dest ), // Templated
		       .reg_pipe0_map9_vc_source(reg_pipe0_map9_vc_source ), // Templated
		       .reg_pipe0_map_en(reg_pipe0_map_en),	 // Templated
		       .reg_pipe0_wr_mode(reg_pipe0_wr_mode[1:0]),
		       .reg_pipe1_drop_ls_le_pkt(reg_pipe1_drop_ls_le_pkt),
		       .reg_pipe1_map0_aggr_id(reg_pipe1_map0_aggr_id), // Templated
		       .reg_pipe1_map0_dt_dest(reg_pipe1_map0_dt_dest ), // Templated
		       .reg_pipe1_map0_dt_source(reg_pipe1_map0_dt_source ), // Templated
		       .reg_pipe1_map0_vc_dest(reg_pipe1_map0_vc_dest ), // Templated
		       .reg_pipe1_map0_vc_source(reg_pipe1_map0_vc_source ), // Templated
		       .reg_pipe1_map10_aggr_id(reg_pipe1_map10_aggr_id), // Templated
		       .reg_pipe1_map10_dt_dest(reg_pipe1_map10_dt_dest), // Templated
		       .reg_pipe1_map10_dt_source(reg_pipe1_map10_dt_source), // Templated
		       .reg_pipe1_map10_vc_dest(reg_pipe1_map10_vc_dest), // Templated
		       .reg_pipe1_map10_vc_source(reg_pipe1_map10_vc_source), // Templated
		       .reg_pipe1_map11_aggr_id(reg_pipe1_map11_aggr_id), // Templated
		       .reg_pipe1_map11_dt_dest(reg_pipe1_map11_dt_dest), // Templated
		       .reg_pipe1_map11_dt_source(reg_pipe1_map11_dt_source), // Templated
		       .reg_pipe1_map11_vc_dest(reg_pipe1_map11_vc_dest), // Templated
		       .reg_pipe1_map11_vc_source(reg_pipe1_map11_vc_source), // Templated
		       .reg_pipe1_map12_aggr_id(reg_pipe1_map12_aggr_id), // Templated
		       .reg_pipe1_map12_dt_dest(reg_pipe1_map12_dt_dest), // Templated
		       .reg_pipe1_map12_dt_source(reg_pipe1_map12_dt_source), // Templated
		       .reg_pipe1_map12_vc_dest(reg_pipe1_map12_vc_dest), // Templated
		       .reg_pipe1_map12_vc_source(reg_pipe1_map12_vc_source), // Templated
		       .reg_pipe1_map13_aggr_id(reg_pipe1_map13_aggr_id), // Templated
		       .reg_pipe1_map13_dt_dest(reg_pipe1_map13_dt_dest), // Templated
		       .reg_pipe1_map13_dt_source(reg_pipe1_map13_dt_source), // Templated
		       .reg_pipe1_map13_vc_dest(reg_pipe1_map13_vc_dest), // Templated
		       .reg_pipe1_map13_vc_source(reg_pipe1_map13_vc_source), // Templated
		       .reg_pipe1_map14_aggr_id(reg_pipe1_map14_aggr_id), // Templated
		       .reg_pipe1_map14_dt_dest(reg_pipe1_map14_dt_dest), // Templated
		       .reg_pipe1_map14_dt_source(reg_pipe1_map14_dt_source), // Templated
		       .reg_pipe1_map14_vc_dest(reg_pipe1_map14_vc_dest), // Templated
		       .reg_pipe1_map14_vc_source(reg_pipe1_map14_vc_source), // Templated
		       .reg_pipe1_map15_aggr_id(reg_pipe1_map15_aggr_id), // Templated
		       .reg_pipe1_map15_dt_dest(reg_pipe1_map15_dt_dest), // Templated
		       .reg_pipe1_map15_dt_source(reg_pipe1_map15_dt_source), // Templated
		       .reg_pipe1_map15_vc_dest(reg_pipe1_map15_vc_dest), // Templated
		       .reg_pipe1_map15_vc_source(reg_pipe1_map15_vc_source), // Templated
		       .reg_pipe1_map1_aggr_id(reg_pipe1_map1_aggr_id), // Templated
		       .reg_pipe1_map1_dt_dest(reg_pipe1_map1_dt_dest ), // Templated
		       .reg_pipe1_map1_dt_source(reg_pipe1_map1_dt_source ), // Templated
		       .reg_pipe1_map1_vc_dest(reg_pipe1_map1_vc_dest ), // Templated
		       .reg_pipe1_map1_vc_source(reg_pipe1_map1_vc_source ), // Templated
		       .reg_pipe1_map2_aggr_id(reg_pipe1_map2_aggr_id), // Templated
		       .reg_pipe1_map2_dt_dest(reg_pipe1_map2_dt_dest ), // Templated
		       .reg_pipe1_map2_dt_source(reg_pipe1_map2_dt_source ), // Templated
		       .reg_pipe1_map2_vc_dest(reg_pipe1_map2_vc_dest ), // Templated
		       .reg_pipe1_map2_vc_source(reg_pipe1_map2_vc_source ), // Templated
		       .reg_pipe1_map3_aggr_id(reg_pipe1_map3_aggr_id), // Templated
		       .reg_pipe1_map3_dt_dest(reg_pipe1_map3_dt_dest ), // Templated
		       .reg_pipe1_map3_dt_source(reg_pipe1_map3_dt_source ), // Templated
		       .reg_pipe1_map3_vc_dest(reg_pipe1_map3_vc_dest ), // Templated
		       .reg_pipe1_map3_vc_source(reg_pipe1_map3_vc_source ), // Templated
		       .reg_pipe1_map4_aggr_id(reg_pipe1_map4_aggr_id), // Templated
		       .reg_pipe1_map4_dt_dest(reg_pipe1_map4_dt_dest ), // Templated
		       .reg_pipe1_map4_dt_source(reg_pipe1_map4_dt_source ), // Templated
		       .reg_pipe1_map4_vc_dest(reg_pipe1_map4_vc_dest ), // Templated
		       .reg_pipe1_map4_vc_source(reg_pipe1_map4_vc_source ), // Templated
		       .reg_pipe1_map5_aggr_id(reg_pipe1_map5_aggr_id), // Templated
		       .reg_pipe1_map5_dt_dest(reg_pipe1_map5_dt_dest ), // Templated
		       .reg_pipe1_map5_dt_source(reg_pipe1_map5_dt_source ), // Templated
		       .reg_pipe1_map5_vc_dest(reg_pipe1_map5_vc_dest ), // Templated
		       .reg_pipe1_map5_vc_source(reg_pipe1_map5_vc_source ), // Templated
		       .reg_pipe1_map6_aggr_id(reg_pipe1_map6_aggr_id), // Templated
		       .reg_pipe1_map6_dt_dest(reg_pipe1_map6_dt_dest ), // Templated
		       .reg_pipe1_map6_dt_source(reg_pipe1_map6_dt_source ), // Templated
		       .reg_pipe1_map6_vc_dest(reg_pipe1_map6_vc_dest ), // Templated
		       .reg_pipe1_map6_vc_source(reg_pipe1_map6_vc_source ), // Templated
		       .reg_pipe1_map7_aggr_id(reg_pipe1_map7_aggr_id), // Templated
		       .reg_pipe1_map7_dt_dest(reg_pipe1_map7_dt_dest ), // Templated
		       .reg_pipe1_map7_dt_source(reg_pipe1_map7_dt_source ), // Templated
		       .reg_pipe1_map7_vc_dest(reg_pipe1_map7_vc_dest ), // Templated
		       .reg_pipe1_map7_vc_source(reg_pipe1_map7_vc_source ), // Templated
		       .reg_pipe1_map8_aggr_id(reg_pipe1_map8_aggr_id), // Templated
		       .reg_pipe1_map8_dt_dest(reg_pipe1_map8_dt_dest ), // Templated
		       .reg_pipe1_map8_dt_source(reg_pipe1_map8_dt_source ), // Templated
		       .reg_pipe1_map8_vc_dest(reg_pipe1_map8_vc_dest ), // Templated
		       .reg_pipe1_map8_vc_source(reg_pipe1_map8_vc_source ), // Templated
		       .reg_pipe1_map9_aggr_id(reg_pipe1_map9_aggr_id), // Templated
		       .reg_pipe1_map9_dt_dest(reg_pipe1_map9_dt_dest ), // Templated
		       .reg_pipe1_map9_dt_source(reg_pipe1_map9_dt_source ), // Templated
		       .reg_pipe1_map9_vc_dest(reg_pipe1_map9_vc_dest ), // Templated
		       .reg_pipe1_map9_vc_source(reg_pipe1_map9_vc_source ), // Templated
		       .reg_pipe1_map_en(reg_pipe1_map_en),	 // Templated
		       .reg_pipe1_wr_mode(reg_pipe1_wr_mode[1:0]),
		       .reg_pipe2_drop_ls_le_pkt(reg_pipe2_drop_ls_le_pkt),
		       .reg_pipe2_map0_aggr_id(reg_pipe2_map0_aggr_id), // Templated
		       .reg_pipe2_map0_dt_dest(reg_pipe2_map0_dt_dest ), // Templated
		       .reg_pipe2_map0_dt_source(reg_pipe2_map0_dt_source ), // Templated
		       .reg_pipe2_map0_vc_dest(reg_pipe2_map0_vc_dest ), // Templated
		       .reg_pipe2_map0_vc_source(reg_pipe2_map0_vc_source ), // Templated
		       .reg_pipe2_map10_aggr_id(reg_pipe2_map10_aggr_id), // Templated
		       .reg_pipe2_map10_dt_dest(reg_pipe2_map10_dt_dest), // Templated
		       .reg_pipe2_map10_dt_source(reg_pipe2_map10_dt_source), // Templated
		       .reg_pipe2_map10_vc_dest(reg_pipe2_map10_vc_dest), // Templated
		       .reg_pipe2_map10_vc_source(reg_pipe2_map10_vc_source), // Templated
		       .reg_pipe2_map11_aggr_id(reg_pipe2_map11_aggr_id), // Templated
		       .reg_pipe2_map11_dt_dest(reg_pipe2_map11_dt_dest), // Templated
		       .reg_pipe2_map11_dt_source(reg_pipe2_map11_dt_source), // Templated
		       .reg_pipe2_map11_vc_dest(reg_pipe2_map11_vc_dest), // Templated
		       .reg_pipe2_map11_vc_source(reg_pipe2_map11_vc_source), // Templated
		       .reg_pipe2_map12_aggr_id(reg_pipe2_map12_aggr_id), // Templated
		       .reg_pipe2_map12_dt_dest(reg_pipe2_map12_dt_dest), // Templated
		       .reg_pipe2_map12_dt_source(reg_pipe2_map12_dt_source), // Templated
		       .reg_pipe2_map12_vc_dest(reg_pipe2_map12_vc_dest), // Templated
		       .reg_pipe2_map12_vc_source(reg_pipe2_map12_vc_source), // Templated
		       .reg_pipe2_map13_aggr_id(reg_pipe2_map13_aggr_id), // Templated
		       .reg_pipe2_map13_dt_dest(reg_pipe2_map13_dt_dest), // Templated
		       .reg_pipe2_map13_dt_source(reg_pipe2_map13_dt_source), // Templated
		       .reg_pipe2_map13_vc_dest(reg_pipe2_map13_vc_dest), // Templated
		       .reg_pipe2_map13_vc_source(reg_pipe2_map13_vc_source), // Templated
		       .reg_pipe2_map14_aggr_id(reg_pipe2_map14_aggr_id), // Templated
		       .reg_pipe2_map14_dt_dest(reg_pipe2_map14_dt_dest), // Templated
		       .reg_pipe2_map14_dt_source(reg_pipe2_map14_dt_source), // Templated
		       .reg_pipe2_map14_vc_dest(reg_pipe2_map14_vc_dest), // Templated
		       .reg_pipe2_map14_vc_source(reg_pipe2_map14_vc_source), // Templated
		       .reg_pipe2_map15_aggr_id(reg_pipe2_map15_aggr_id), // Templated
		       .reg_pipe2_map15_dt_dest(reg_pipe2_map15_dt_dest), // Templated
		       .reg_pipe2_map15_dt_source(reg_pipe2_map15_dt_source), // Templated
		       .reg_pipe2_map15_vc_dest(reg_pipe2_map15_vc_dest), // Templated
		       .reg_pipe2_map15_vc_source(reg_pipe2_map15_vc_source), // Templated
		       .reg_pipe2_map1_aggr_id(reg_pipe2_map1_aggr_id), // Templated
		       .reg_pipe2_map1_dt_dest(reg_pipe2_map1_dt_dest ), // Templated
		       .reg_pipe2_map1_dt_source(reg_pipe2_map1_dt_source ), // Templated
		       .reg_pipe2_map1_vc_dest(reg_pipe2_map1_vc_dest ), // Templated
		       .reg_pipe2_map1_vc_source(reg_pipe2_map1_vc_source ), // Templated
		       .reg_pipe2_map2_aggr_id(reg_pipe2_map2_aggr_id), // Templated
		       .reg_pipe2_map2_dt_dest(reg_pipe2_map2_dt_dest ), // Templated
		       .reg_pipe2_map2_dt_source(reg_pipe2_map2_dt_source ), // Templated
		       .reg_pipe2_map2_vc_dest(reg_pipe2_map2_vc_dest ), // Templated
		       .reg_pipe2_map2_vc_source(reg_pipe2_map2_vc_source ), // Templated
		       .reg_pipe2_map3_aggr_id(reg_pipe2_map3_aggr_id), // Templated
		       .reg_pipe2_map3_dt_dest(reg_pipe2_map3_dt_dest ), // Templated
		       .reg_pipe2_map3_dt_source(reg_pipe2_map3_dt_source ), // Templated
		       .reg_pipe2_map3_vc_dest(reg_pipe2_map3_vc_dest ), // Templated
		       .reg_pipe2_map3_vc_source(reg_pipe2_map3_vc_source ), // Templated
		       .reg_pipe2_map4_aggr_id(reg_pipe2_map4_aggr_id), // Templated
		       .reg_pipe2_map4_dt_dest(reg_pipe2_map4_dt_dest ), // Templated
		       .reg_pipe2_map4_dt_source(reg_pipe2_map4_dt_source ), // Templated
		       .reg_pipe2_map4_vc_dest(reg_pipe2_map4_vc_dest ), // Templated
		       .reg_pipe2_map4_vc_source(reg_pipe2_map4_vc_source ), // Templated
		       .reg_pipe2_map5_aggr_id(reg_pipe2_map5_aggr_id), // Templated
		       .reg_pipe2_map5_dt_dest(reg_pipe2_map5_dt_dest ), // Templated
		       .reg_pipe2_map5_dt_source(reg_pipe2_map5_dt_source ), // Templated
		       .reg_pipe2_map5_vc_dest(reg_pipe2_map5_vc_dest ), // Templated
		       .reg_pipe2_map5_vc_source(reg_pipe2_map5_vc_source ), // Templated
		       .reg_pipe2_map6_aggr_id(reg_pipe2_map6_aggr_id), // Templated
		       .reg_pipe2_map6_dt_dest(reg_pipe2_map6_dt_dest ), // Templated
		       .reg_pipe2_map6_dt_source(reg_pipe2_map6_dt_source ), // Templated
		       .reg_pipe2_map6_vc_dest(reg_pipe2_map6_vc_dest ), // Templated
		       .reg_pipe2_map6_vc_source(reg_pipe2_map6_vc_source ), // Templated
		       .reg_pipe2_map7_aggr_id(reg_pipe2_map7_aggr_id), // Templated
		       .reg_pipe2_map7_dt_dest(reg_pipe2_map7_dt_dest ), // Templated
		       .reg_pipe2_map7_dt_source(reg_pipe2_map7_dt_source ), // Templated
		       .reg_pipe2_map7_vc_dest(reg_pipe2_map7_vc_dest ), // Templated
		       .reg_pipe2_map7_vc_source(reg_pipe2_map7_vc_source ), // Templated
		       .reg_pipe2_map8_aggr_id(reg_pipe2_map8_aggr_id), // Templated
		       .reg_pipe2_map8_dt_dest(reg_pipe2_map8_dt_dest ), // Templated
		       .reg_pipe2_map8_dt_source(reg_pipe2_map8_dt_source ), // Templated
		       .reg_pipe2_map8_vc_dest(reg_pipe2_map8_vc_dest ), // Templated
		       .reg_pipe2_map8_vc_source(reg_pipe2_map8_vc_source ), // Templated
		       .reg_pipe2_map9_aggr_id(reg_pipe2_map9_aggr_id), // Templated
		       .reg_pipe2_map9_dt_dest(reg_pipe2_map9_dt_dest ), // Templated
		       .reg_pipe2_map9_dt_source(reg_pipe2_map9_dt_source ), // Templated
		       .reg_pipe2_map9_vc_dest(reg_pipe2_map9_vc_dest ), // Templated
		       .reg_pipe2_map9_vc_source(reg_pipe2_map9_vc_source ), // Templated
		       .reg_pipe2_map_en(reg_pipe2_map_en),	 // Templated
		       .reg_pipe2_wr_mode(reg_pipe2_wr_mode[1:0]),
		       .reg_pipe3_drop_ls_le_pkt(reg_pipe3_drop_ls_le_pkt),
		       .reg_pipe3_map0_aggr_id(reg_pipe3_map0_aggr_id), // Templated
		       .reg_pipe3_map0_dt_dest(reg_pipe3_map0_dt_dest ), // Templated
		       .reg_pipe3_map0_dt_source(reg_pipe3_map0_dt_source ), // Templated
		       .reg_pipe3_map0_vc_dest(reg_pipe3_map0_vc_dest ), // Templated
		       .reg_pipe3_map0_vc_source(reg_pipe3_map0_vc_source ), // Templated
		       .reg_pipe3_map10_aggr_id(reg_pipe3_map10_aggr_id), // Templated
		       .reg_pipe3_map10_dt_dest(reg_pipe3_map10_dt_dest), // Templated
		       .reg_pipe3_map10_dt_source(reg_pipe3_map10_dt_source), // Templated
		       .reg_pipe3_map10_vc_dest(reg_pipe3_map10_vc_dest), // Templated
		       .reg_pipe3_map10_vc_source(reg_pipe3_map10_vc_source), // Templated
		       .reg_pipe3_map11_aggr_id(reg_pipe3_map11_aggr_id), // Templated
		       .reg_pipe3_map11_dt_dest(reg_pipe3_map11_dt_dest), // Templated
		       .reg_pipe3_map11_dt_source(reg_pipe3_map11_dt_source), // Templated
		       .reg_pipe3_map11_vc_dest(reg_pipe3_map11_vc_dest), // Templated
		       .reg_pipe3_map11_vc_source(reg_pipe3_map11_vc_source), // Templated
		       .reg_pipe3_map12_aggr_id(reg_pipe3_map12_aggr_id), // Templated
		       .reg_pipe3_map12_dt_dest(reg_pipe3_map12_dt_dest), // Templated
		       .reg_pipe3_map12_dt_source(reg_pipe3_map12_dt_source), // Templated
		       .reg_pipe3_map12_vc_dest(reg_pipe3_map12_vc_dest), // Templated
		       .reg_pipe3_map12_vc_source(reg_pipe3_map12_vc_source), // Templated
		       .reg_pipe3_map13_aggr_id(reg_pipe3_map13_aggr_id), // Templated
		       .reg_pipe3_map13_dt_dest(reg_pipe3_map13_dt_dest), // Templated
		       .reg_pipe3_map13_dt_source(reg_pipe3_map13_dt_source), // Templated
		       .reg_pipe3_map13_vc_dest(reg_pipe3_map13_vc_dest), // Templated
		       .reg_pipe3_map13_vc_source(reg_pipe3_map13_vc_source), // Templated
		       .reg_pipe3_map14_aggr_id(reg_pipe3_map14_aggr_id), // Templated
		       .reg_pipe3_map14_dt_dest(reg_pipe3_map14_dt_dest), // Templated
		       .reg_pipe3_map14_dt_source(reg_pipe3_map14_dt_source), // Templated
		       .reg_pipe3_map14_vc_dest(reg_pipe3_map14_vc_dest), // Templated
		       .reg_pipe3_map14_vc_source(reg_pipe3_map14_vc_source), // Templated
		       .reg_pipe3_map15_aggr_id(reg_pipe3_map15_aggr_id), // Templated
		       .reg_pipe3_map15_dt_dest(reg_pipe3_map15_dt_dest), // Templated
		       .reg_pipe3_map15_dt_source(reg_pipe3_map15_dt_source), // Templated
		       .reg_pipe3_map15_vc_dest(reg_pipe3_map15_vc_dest), // Templated
		       .reg_pipe3_map15_vc_source(reg_pipe3_map15_vc_source), // Templated
		       .reg_pipe3_map1_aggr_id(reg_pipe3_map1_aggr_id), // Templated
		       .reg_pipe3_map1_dt_dest(reg_pipe3_map1_dt_dest ), // Templated
		       .reg_pipe3_map1_dt_source(reg_pipe3_map1_dt_source ), // Templated
		       .reg_pipe3_map1_vc_dest(reg_pipe3_map1_vc_dest ), // Templated
		       .reg_pipe3_map1_vc_source(reg_pipe3_map1_vc_source ), // Templated
		       .reg_pipe3_map2_aggr_id(reg_pipe3_map2_aggr_id), // Templated
		       .reg_pipe3_map2_dt_dest(reg_pipe3_map2_dt_dest ), // Templated
		       .reg_pipe3_map2_dt_source(reg_pipe3_map2_dt_source ), // Templated
		       .reg_pipe3_map2_vc_dest(reg_pipe3_map2_vc_dest ), // Templated
		       .reg_pipe3_map2_vc_source(reg_pipe3_map2_vc_source ), // Templated
		       .reg_pipe3_map3_aggr_id(reg_pipe3_map3_aggr_id), // Templated
		       .reg_pipe3_map3_dt_dest(reg_pipe3_map3_dt_dest ), // Templated
		       .reg_pipe3_map3_dt_source(reg_pipe3_map3_dt_source ), // Templated
		       .reg_pipe3_map3_vc_dest(reg_pipe3_map3_vc_dest ), // Templated
		       .reg_pipe3_map3_vc_source(reg_pipe3_map3_vc_source ), // Templated
		       .reg_pipe3_map4_aggr_id(reg_pipe3_map4_aggr_id), // Templated
		       .reg_pipe3_map4_dt_dest(reg_pipe3_map4_dt_dest ), // Templated
		       .reg_pipe3_map4_dt_source(reg_pipe3_map4_dt_source ), // Templated
		       .reg_pipe3_map4_vc_dest(reg_pipe3_map4_vc_dest ), // Templated
		       .reg_pipe3_map4_vc_source(reg_pipe3_map4_vc_source ), // Templated
		       .reg_pipe3_map5_aggr_id(reg_pipe3_map5_aggr_id), // Templated
		       .reg_pipe3_map5_dt_dest(reg_pipe3_map5_dt_dest ), // Templated
		       .reg_pipe3_map5_dt_source(reg_pipe3_map5_dt_source ), // Templated
		       .reg_pipe3_map5_vc_dest(reg_pipe3_map5_vc_dest ), // Templated
		       .reg_pipe3_map5_vc_source(reg_pipe3_map5_vc_source ), // Templated
		       .reg_pipe3_map6_aggr_id(reg_pipe3_map6_aggr_id), // Templated
		       .reg_pipe3_map6_dt_dest(reg_pipe3_map6_dt_dest ), // Templated
		       .reg_pipe3_map6_dt_source(reg_pipe3_map6_dt_source ), // Templated
		       .reg_pipe3_map6_vc_dest(reg_pipe3_map6_vc_dest ), // Templated
		       .reg_pipe3_map6_vc_source(reg_pipe3_map6_vc_source ), // Templated
		       .reg_pipe3_map7_aggr_id(reg_pipe3_map7_aggr_id), // Templated
		       .reg_pipe3_map7_dt_dest(reg_pipe3_map7_dt_dest ), // Templated
		       .reg_pipe3_map7_dt_source(reg_pipe3_map7_dt_source ), // Templated
		       .reg_pipe3_map7_vc_dest(reg_pipe3_map7_vc_dest ), // Templated
		       .reg_pipe3_map7_vc_source(reg_pipe3_map7_vc_source ), // Templated
		       .reg_pipe3_map8_aggr_id(reg_pipe3_map8_aggr_id), // Templated
		       .reg_pipe3_map8_dt_dest(reg_pipe3_map8_dt_dest ), // Templated
		       .reg_pipe3_map8_dt_source(reg_pipe3_map8_dt_source ), // Templated
		       .reg_pipe3_map8_vc_dest(reg_pipe3_map8_vc_dest ), // Templated
		       .reg_pipe3_map8_vc_source(reg_pipe3_map8_vc_source ), // Templated
		       .reg_pipe3_map9_aggr_id(reg_pipe3_map9_aggr_id), // Templated
		       .reg_pipe3_map9_dt_dest(reg_pipe3_map9_dt_dest ), // Templated
		       .reg_pipe3_map9_dt_source(reg_pipe3_map9_dt_source ), // Templated
		       .reg_pipe3_map9_vc_dest(reg_pipe3_map9_vc_dest ), // Templated
		       .reg_pipe3_map9_vc_source(reg_pipe3_map9_vc_source ), // Templated
		       .reg_pipe3_map_en(reg_pipe3_map_en),	 // Templated
		       .reg_pipe3_wr_mode(reg_pipe3_wr_mode[1:0]),
		       .reg_pipe4_drop_ls_le_pkt(reg_pipe4_drop_ls_le_pkt),
		       .reg_pipe4_map0_aggr_id(reg_pipe4_map0_aggr_id[3:0]),
		       .reg_pipe4_map0_dt_dest(reg_pipe4_map0_dt_dest ), // Templated
		       .reg_pipe4_map0_dt_source(reg_pipe4_map0_dt_source ), // Templated
		       .reg_pipe4_map0_vc_dest(reg_pipe4_map0_vc_dest ), // Templated
		       .reg_pipe4_map0_vc_source(reg_pipe4_map0_vc_source ), // Templated
		       .reg_pipe4_map10_aggr_id(reg_pipe4_map10_aggr_id[3:0]),
		       .reg_pipe4_map10_dt_dest(reg_pipe4_map10_dt_dest), // Templated
		       .reg_pipe4_map10_dt_source(reg_pipe4_map10_dt_source), // Templated
		       .reg_pipe4_map10_vc_dest(reg_pipe4_map10_vc_dest), // Templated
		       .reg_pipe4_map10_vc_source(reg_pipe4_map10_vc_source), // Templated
		       .reg_pipe4_map11_aggr_id(reg_pipe4_map11_aggr_id[3:0]),
		       .reg_pipe4_map11_dt_dest(reg_pipe4_map11_dt_dest), // Templated
		       .reg_pipe4_map11_dt_source(reg_pipe4_map11_dt_source), // Templated
		       .reg_pipe4_map11_vc_dest(reg_pipe4_map11_vc_dest), // Templated
		       .reg_pipe4_map11_vc_source(reg_pipe4_map11_vc_source), // Templated
		       .reg_pipe4_map12_aggr_id(reg_pipe4_map12_aggr_id[3:0]),
		       .reg_pipe4_map12_dt_dest(reg_pipe4_map12_dt_dest), // Templated
		       .reg_pipe4_map12_dt_source(reg_pipe4_map12_dt_source), // Templated
		       .reg_pipe4_map12_vc_dest(reg_pipe4_map12_vc_dest), // Templated
		       .reg_pipe4_map12_vc_source(reg_pipe4_map12_vc_source), // Templated
		       .reg_pipe4_map13_aggr_id(reg_pipe4_map13_aggr_id[3:0]),
		       .reg_pipe4_map13_dt_dest(reg_pipe4_map13_dt_dest), // Templated
		       .reg_pipe4_map13_dt_source(reg_pipe4_map13_dt_source), // Templated
		       .reg_pipe4_map13_vc_dest(reg_pipe4_map13_vc_dest), // Templated
		       .reg_pipe4_map13_vc_source(reg_pipe4_map13_vc_source), // Templated
		       .reg_pipe4_map14_aggr_id(reg_pipe4_map14_aggr_id[3:0]),
		       .reg_pipe4_map14_dt_dest(reg_pipe4_map14_dt_dest), // Templated
		       .reg_pipe4_map14_dt_source(reg_pipe4_map14_dt_source), // Templated
		       .reg_pipe4_map14_vc_dest(reg_pipe4_map14_vc_dest), // Templated
		       .reg_pipe4_map14_vc_source(reg_pipe4_map14_vc_source), // Templated
		       .reg_pipe4_map15_aggr_id(reg_pipe4_map15_aggr_id[3:0]),
		       .reg_pipe4_map15_dt_dest(reg_pipe4_map15_dt_dest), // Templated
		       .reg_pipe4_map15_dt_source(reg_pipe4_map15_dt_source), // Templated
		       .reg_pipe4_map15_vc_dest(reg_pipe4_map15_vc_dest), // Templated
		       .reg_pipe4_map15_vc_source(reg_pipe4_map15_vc_source), // Templated
		       .reg_pipe4_map1_aggr_id(reg_pipe4_map1_aggr_id[3:0]),
		       .reg_pipe4_map1_dt_dest(reg_pipe4_map1_dt_dest ), // Templated
		       .reg_pipe4_map1_dt_source(reg_pipe4_map1_dt_source ), // Templated
		       .reg_pipe4_map1_vc_dest(reg_pipe4_map1_vc_dest ), // Templated
		       .reg_pipe4_map1_vc_source(reg_pipe4_map1_vc_source ), // Templated
		       .reg_pipe4_map2_aggr_id(reg_pipe4_map2_aggr_id[3:0]),
		       .reg_pipe4_map2_dt_dest(reg_pipe4_map2_dt_dest ), // Templated
		       .reg_pipe4_map2_dt_source(reg_pipe4_map2_dt_source ), // Templated
		       .reg_pipe4_map2_vc_dest(reg_pipe4_map2_vc_dest ), // Templated
		       .reg_pipe4_map2_vc_source(reg_pipe4_map2_vc_source ), // Templated
		       .reg_pipe4_map3_aggr_id(reg_pipe4_map3_aggr_id[3:0]),
		       .reg_pipe4_map3_dt_dest(reg_pipe4_map3_dt_dest ), // Templated
		       .reg_pipe4_map3_dt_source(reg_pipe4_map3_dt_source ), // Templated
		       .reg_pipe4_map3_vc_dest(reg_pipe4_map3_vc_dest ), // Templated
		       .reg_pipe4_map3_vc_source(reg_pipe4_map3_vc_source ), // Templated
		       .reg_pipe4_map4_aggr_id(reg_pipe4_map4_aggr_id[3:0]),
		       .reg_pipe4_map4_dt_dest(reg_pipe4_map4_dt_dest ), // Templated
		       .reg_pipe4_map4_dt_source(reg_pipe4_map4_dt_source ), // Templated
		       .reg_pipe4_map4_vc_dest(reg_pipe4_map4_vc_dest ), // Templated
		       .reg_pipe4_map4_vc_source(reg_pipe4_map4_vc_source ), // Templated
		       .reg_pipe4_map5_aggr_id(reg_pipe4_map5_aggr_id[3:0]),
		       .reg_pipe4_map5_dt_dest(reg_pipe4_map5_dt_dest ), // Templated
		       .reg_pipe4_map5_dt_source(reg_pipe4_map5_dt_source ), // Templated
		       .reg_pipe4_map5_vc_dest(reg_pipe4_map5_vc_dest ), // Templated
		       .reg_pipe4_map5_vc_source(reg_pipe4_map5_vc_source ), // Templated
		       .reg_pipe4_map6_aggr_id(reg_pipe4_map6_aggr_id[3:0]),
		       .reg_pipe4_map6_dt_dest(reg_pipe4_map6_dt_dest ), // Templated
		       .reg_pipe4_map6_dt_source(reg_pipe4_map6_dt_source ), // Templated
		       .reg_pipe4_map6_vc_dest(reg_pipe4_map6_vc_dest ), // Templated
		       .reg_pipe4_map6_vc_source(reg_pipe4_map6_vc_source ), // Templated
		       .reg_pipe4_map7_aggr_id(reg_pipe4_map7_aggr_id[3:0]),
		       .reg_pipe4_map7_dt_dest(reg_pipe4_map7_dt_dest ), // Templated
		       .reg_pipe4_map7_dt_source(reg_pipe4_map7_dt_source ), // Templated
		       .reg_pipe4_map7_vc_dest(reg_pipe4_map7_vc_dest ), // Templated
		       .reg_pipe4_map7_vc_source(reg_pipe4_map7_vc_source ), // Templated
		       .reg_pipe4_map8_aggr_id(reg_pipe4_map8_aggr_id[3:0]),
		       .reg_pipe4_map8_dt_dest(reg_pipe4_map8_dt_dest ), // Templated
		       .reg_pipe4_map8_dt_source(reg_pipe4_map8_dt_source ), // Templated
		       .reg_pipe4_map8_vc_dest(reg_pipe4_map8_vc_dest ), // Templated
		       .reg_pipe4_map8_vc_source(reg_pipe4_map8_vc_source ), // Templated
		       .reg_pipe4_map9_aggr_id(reg_pipe4_map9_aggr_id[3:0]),
		       .reg_pipe4_map9_dt_dest(reg_pipe4_map9_dt_dest ), // Templated
		       .reg_pipe4_map9_dt_source(reg_pipe4_map9_dt_source ), // Templated
		       .reg_pipe4_map9_vc_dest(reg_pipe4_map9_vc_dest ), // Templated
		       .reg_pipe4_map9_vc_source(reg_pipe4_map9_vc_source ), // Templated
		       .reg_pipe4_map_en(reg_pipe4_map_en),	 // Templated
		       .reg_pipe4_wr_mode(reg_pipe4_wr_mode[1:0]),
		       .reg_pipe5_drop_ls_le_pkt(reg_pipe5_drop_ls_le_pkt),
		       .reg_pipe5_map0_aggr_id(reg_pipe5_map0_aggr_id[3:0]),
		       .reg_pipe5_map0_dt_dest(reg_pipe5_map0_dt_dest ), // Templated
		       .reg_pipe5_map0_dt_source(reg_pipe5_map0_dt_source ), // Templated
		       .reg_pipe5_map0_vc_dest(reg_pipe5_map0_vc_dest ), // Templated
		       .reg_pipe5_map0_vc_source(reg_pipe5_map0_vc_source ), // Templated
		       .reg_pipe5_map10_aggr_id(reg_pipe5_map10_aggr_id[3:0]),
		       .reg_pipe5_map10_dt_dest(reg_pipe5_map10_dt_dest), // Templated
		       .reg_pipe5_map10_dt_source(reg_pipe5_map10_dt_source), // Templated
		       .reg_pipe5_map10_vc_dest(reg_pipe5_map10_vc_dest), // Templated
		       .reg_pipe5_map10_vc_source(reg_pipe5_map10_vc_source), // Templated
		       .reg_pipe5_map11_aggr_id(reg_pipe5_map11_aggr_id[3:0]),
		       .reg_pipe5_map11_dt_dest(reg_pipe5_map11_dt_dest), // Templated
		       .reg_pipe5_map11_dt_source(reg_pipe5_map11_dt_source), // Templated
		       .reg_pipe5_map11_vc_dest(reg_pipe5_map11_vc_dest), // Templated
		       .reg_pipe5_map11_vc_source(reg_pipe5_map11_vc_source), // Templated
		       .reg_pipe5_map12_aggr_id(reg_pipe5_map12_aggr_id[3:0]),
		       .reg_pipe5_map12_dt_dest(reg_pipe5_map12_dt_dest), // Templated
		       .reg_pipe5_map12_dt_source(reg_pipe5_map12_dt_source), // Templated
		       .reg_pipe5_map12_vc_dest(reg_pipe5_map12_vc_dest), // Templated
		       .reg_pipe5_map12_vc_source(reg_pipe5_map12_vc_source), // Templated
		       .reg_pipe5_map13_aggr_id(reg_pipe5_map13_aggr_id[3:0]),
		       .reg_pipe5_map13_dt_dest(reg_pipe5_map13_dt_dest), // Templated
		       .reg_pipe5_map13_dt_source(reg_pipe5_map13_dt_source), // Templated
		       .reg_pipe5_map13_vc_dest(reg_pipe5_map13_vc_dest), // Templated
		       .reg_pipe5_map13_vc_source(reg_pipe5_map13_vc_source), // Templated
		       .reg_pipe5_map14_aggr_id(reg_pipe5_map14_aggr_id[3:0]),
		       .reg_pipe5_map14_dt_dest(reg_pipe5_map14_dt_dest), // Templated
		       .reg_pipe5_map14_dt_source(reg_pipe5_map14_dt_source), // Templated
		       .reg_pipe5_map14_vc_dest(reg_pipe5_map14_vc_dest), // Templated
		       .reg_pipe5_map14_vc_source(reg_pipe5_map14_vc_source), // Templated
		       .reg_pipe5_map15_aggr_id(reg_pipe5_map15_aggr_id[3:0]),
		       .reg_pipe5_map15_dt_dest(reg_pipe5_map15_dt_dest), // Templated
		       .reg_pipe5_map15_dt_source(reg_pipe5_map15_dt_source), // Templated
		       .reg_pipe5_map15_vc_dest(reg_pipe5_map15_vc_dest), // Templated
		       .reg_pipe5_map15_vc_source(reg_pipe5_map15_vc_source), // Templated
		       .reg_pipe5_map1_aggr_id(reg_pipe5_map1_aggr_id[3:0]),
		       .reg_pipe5_map1_dt_dest(reg_pipe5_map1_dt_dest ), // Templated
		       .reg_pipe5_map1_dt_source(reg_pipe5_map1_dt_source ), // Templated
		       .reg_pipe5_map1_vc_dest(reg_pipe5_map1_vc_dest ), // Templated
		       .reg_pipe5_map1_vc_source(reg_pipe5_map1_vc_source ), // Templated
		       .reg_pipe5_map2_aggr_id(reg_pipe5_map2_aggr_id[3:0]),
		       .reg_pipe5_map2_dt_dest(reg_pipe5_map2_dt_dest ), // Templated
		       .reg_pipe5_map2_dt_source(reg_pipe5_map2_dt_source ), // Templated
		       .reg_pipe5_map2_vc_dest(reg_pipe5_map2_vc_dest ), // Templated
		       .reg_pipe5_map2_vc_source(reg_pipe5_map2_vc_source ), // Templated
		       .reg_pipe5_map3_aggr_id(reg_pipe5_map3_aggr_id[3:0]),
		       .reg_pipe5_map3_dt_dest(reg_pipe5_map3_dt_dest ), // Templated
		       .reg_pipe5_map3_dt_source(reg_pipe5_map3_dt_source ), // Templated
		       .reg_pipe5_map3_vc_dest(reg_pipe5_map3_vc_dest ), // Templated
		       .reg_pipe5_map3_vc_source(reg_pipe5_map3_vc_source ), // Templated
		       .reg_pipe5_map4_aggr_id(reg_pipe5_map4_aggr_id[3:0]),
		       .reg_pipe5_map4_dt_dest(reg_pipe5_map4_dt_dest ), // Templated
		       .reg_pipe5_map4_dt_source(reg_pipe5_map4_dt_source ), // Templated
		       .reg_pipe5_map4_vc_dest(reg_pipe5_map4_vc_dest ), // Templated
		       .reg_pipe5_map4_vc_source(reg_pipe5_map4_vc_source ), // Templated
		       .reg_pipe5_map5_aggr_id(reg_pipe5_map5_aggr_id[3:0]),
		       .reg_pipe5_map5_dt_dest(reg_pipe5_map5_dt_dest ), // Templated
		       .reg_pipe5_map5_dt_source(reg_pipe5_map5_dt_source ), // Templated
		       .reg_pipe5_map5_vc_dest(reg_pipe5_map5_vc_dest ), // Templated
		       .reg_pipe5_map5_vc_source(reg_pipe5_map5_vc_source ), // Templated
		       .reg_pipe5_map6_aggr_id(reg_pipe5_map6_aggr_id[3:0]),
		       .reg_pipe5_map6_dt_dest(reg_pipe5_map6_dt_dest ), // Templated
		       .reg_pipe5_map6_dt_source(reg_pipe5_map6_dt_source ), // Templated
		       .reg_pipe5_map6_vc_dest(reg_pipe5_map6_vc_dest ), // Templated
		       .reg_pipe5_map6_vc_source(reg_pipe5_map6_vc_source ), // Templated
		       .reg_pipe5_map7_aggr_id(reg_pipe5_map7_aggr_id[3:0]),
		       .reg_pipe5_map7_dt_dest(reg_pipe5_map7_dt_dest ), // Templated
		       .reg_pipe5_map7_dt_source(reg_pipe5_map7_dt_source ), // Templated
		       .reg_pipe5_map7_vc_dest(reg_pipe5_map7_vc_dest ), // Templated
		       .reg_pipe5_map7_vc_source(reg_pipe5_map7_vc_source ), // Templated
		       .reg_pipe5_map8_aggr_id(reg_pipe5_map8_aggr_id[3:0]),
		       .reg_pipe5_map8_dt_dest(reg_pipe5_map8_dt_dest ), // Templated
		       .reg_pipe5_map8_dt_source(reg_pipe5_map8_dt_source ), // Templated
		       .reg_pipe5_map8_vc_dest(reg_pipe5_map8_vc_dest ), // Templated
		       .reg_pipe5_map8_vc_source(reg_pipe5_map8_vc_source ), // Templated
		       .reg_pipe5_map9_aggr_id(reg_pipe5_map9_aggr_id[3:0]),
		       .reg_pipe5_map9_dt_dest(reg_pipe5_map9_dt_dest ), // Templated
		       .reg_pipe5_map9_dt_source(reg_pipe5_map9_dt_source ), // Templated
		       .reg_pipe5_map9_vc_dest(reg_pipe5_map9_vc_dest ), // Templated
		       .reg_pipe5_map9_vc_source(reg_pipe5_map9_vc_source ), // Templated
		       .reg_pipe5_map_en(reg_pipe5_map_en),	 // Templated
		       .reg_pipe5_wr_mode(reg_pipe5_wr_mode[1:0]),
		       .reg_pipe6_drop_ls_le_pkt(reg_pipe6_drop_ls_le_pkt),
		       .reg_pipe6_map0_aggr_id(reg_pipe6_map0_aggr_id[3:0]),
		       .reg_pipe6_map0_dt_dest(reg_pipe6_map0_dt_dest ), // Templated
		       .reg_pipe6_map0_dt_source(reg_pipe6_map0_dt_source ), // Templated
		       .reg_pipe6_map0_vc_dest(reg_pipe6_map0_vc_dest ), // Templated
		       .reg_pipe6_map0_vc_source(reg_pipe6_map0_vc_source ), // Templated
		       .reg_pipe6_map10_aggr_id(reg_pipe6_map10_aggr_id[3:0]),
		       .reg_pipe6_map10_dt_dest(reg_pipe6_map10_dt_dest), // Templated
		       .reg_pipe6_map10_dt_source(reg_pipe6_map10_dt_source), // Templated
		       .reg_pipe6_map10_vc_dest(reg_pipe6_map10_vc_dest), // Templated
		       .reg_pipe6_map10_vc_source(reg_pipe6_map10_vc_source), // Templated
		       .reg_pipe6_map11_aggr_id(reg_pipe6_map11_aggr_id[3:0]),
		       .reg_pipe6_map11_dt_dest(reg_pipe6_map11_dt_dest), // Templated
		       .reg_pipe6_map11_dt_source(reg_pipe6_map11_dt_source), // Templated
		       .reg_pipe6_map11_vc_dest(reg_pipe6_map11_vc_dest), // Templated
		       .reg_pipe6_map11_vc_source(reg_pipe6_map11_vc_source), // Templated
		       .reg_pipe6_map12_aggr_id(reg_pipe6_map12_aggr_id[3:0]),
		       .reg_pipe6_map12_dt_dest(reg_pipe6_map12_dt_dest), // Templated
		       .reg_pipe6_map12_dt_source(reg_pipe6_map12_dt_source), // Templated
		       .reg_pipe6_map12_vc_dest(reg_pipe6_map12_vc_dest), // Templated
		       .reg_pipe6_map12_vc_source(reg_pipe6_map12_vc_source), // Templated
		       .reg_pipe6_map13_aggr_id(reg_pipe6_map13_aggr_id[3:0]),
		       .reg_pipe6_map13_dt_dest(reg_pipe6_map13_dt_dest), // Templated
		       .reg_pipe6_map13_dt_source(reg_pipe6_map13_dt_source), // Templated
		       .reg_pipe6_map13_vc_dest(reg_pipe6_map13_vc_dest), // Templated
		       .reg_pipe6_map13_vc_source(reg_pipe6_map13_vc_source), // Templated
		       .reg_pipe6_map14_aggr_id(reg_pipe6_map14_aggr_id[3:0]),
		       .reg_pipe6_map14_dt_dest(reg_pipe6_map14_dt_dest), // Templated
		       .reg_pipe6_map14_dt_source(reg_pipe6_map14_dt_source), // Templated
		       .reg_pipe6_map14_vc_dest(reg_pipe6_map14_vc_dest), // Templated
		       .reg_pipe6_map14_vc_source(reg_pipe6_map14_vc_source), // Templated
		       .reg_pipe6_map15_aggr_id(reg_pipe6_map15_aggr_id[3:0]),
		       .reg_pipe6_map15_dt_dest(reg_pipe6_map15_dt_dest), // Templated
		       .reg_pipe6_map15_dt_source(reg_pipe6_map15_dt_source), // Templated
		       .reg_pipe6_map15_vc_dest(reg_pipe6_map15_vc_dest), // Templated
		       .reg_pipe6_map15_vc_source(reg_pipe6_map15_vc_source), // Templated
		       .reg_pipe6_map1_aggr_id(reg_pipe6_map1_aggr_id[3:0]),
		       .reg_pipe6_map1_dt_dest(reg_pipe6_map1_dt_dest ), // Templated
		       .reg_pipe6_map1_dt_source(reg_pipe6_map1_dt_source ), // Templated
		       .reg_pipe6_map1_vc_dest(reg_pipe6_map1_vc_dest ), // Templated
		       .reg_pipe6_map1_vc_source(reg_pipe6_map1_vc_source ), // Templated
		       .reg_pipe6_map2_aggr_id(reg_pipe6_map2_aggr_id[3:0]),
		       .reg_pipe6_map2_dt_dest(reg_pipe6_map2_dt_dest ), // Templated
		       .reg_pipe6_map2_dt_source(reg_pipe6_map2_dt_source ), // Templated
		       .reg_pipe6_map2_vc_dest(reg_pipe6_map2_vc_dest ), // Templated
		       .reg_pipe6_map2_vc_source(reg_pipe6_map2_vc_source ), // Templated
		       .reg_pipe6_map3_aggr_id(reg_pipe6_map3_aggr_id[3:0]),
		       .reg_pipe6_map3_dt_dest(reg_pipe6_map3_dt_dest ), // Templated
		       .reg_pipe6_map3_dt_source(reg_pipe6_map3_dt_source ), // Templated
		       .reg_pipe6_map3_vc_dest(reg_pipe6_map3_vc_dest ), // Templated
		       .reg_pipe6_map3_vc_source(reg_pipe6_map3_vc_source ), // Templated
		       .reg_pipe6_map4_aggr_id(reg_pipe6_map4_aggr_id[3:0]),
		       .reg_pipe6_map4_dt_dest(reg_pipe6_map4_dt_dest ), // Templated
		       .reg_pipe6_map4_dt_source(reg_pipe6_map4_dt_source ), // Templated
		       .reg_pipe6_map4_vc_dest(reg_pipe6_map4_vc_dest ), // Templated
		       .reg_pipe6_map4_vc_source(reg_pipe6_map4_vc_source ), // Templated
		       .reg_pipe6_map5_aggr_id(reg_pipe6_map5_aggr_id[3:0]),
		       .reg_pipe6_map5_dt_dest(reg_pipe6_map5_dt_dest ), // Templated
		       .reg_pipe6_map5_dt_source(reg_pipe6_map5_dt_source ), // Templated
		       .reg_pipe6_map5_vc_dest(reg_pipe6_map5_vc_dest ), // Templated
		       .reg_pipe6_map5_vc_source(reg_pipe6_map5_vc_source ), // Templated
		       .reg_pipe6_map6_aggr_id(reg_pipe6_map6_aggr_id[3:0]),
		       .reg_pipe6_map6_dt_dest(reg_pipe6_map6_dt_dest ), // Templated
		       .reg_pipe6_map6_dt_source(reg_pipe6_map6_dt_source ), // Templated
		       .reg_pipe6_map6_vc_dest(reg_pipe6_map6_vc_dest ), // Templated
		       .reg_pipe6_map6_vc_source(reg_pipe6_map6_vc_source ), // Templated
		       .reg_pipe6_map7_aggr_id(reg_pipe6_map7_aggr_id[3:0]),
		       .reg_pipe6_map7_dt_dest(reg_pipe6_map7_dt_dest ), // Templated
		       .reg_pipe6_map7_dt_source(reg_pipe6_map7_dt_source ), // Templated
		       .reg_pipe6_map7_vc_dest(reg_pipe6_map7_vc_dest ), // Templated
		       .reg_pipe6_map7_vc_source(reg_pipe6_map7_vc_source ), // Templated
		       .reg_pipe6_map8_aggr_id(reg_pipe6_map8_aggr_id[3:0]),
		       .reg_pipe6_map8_dt_dest(reg_pipe6_map8_dt_dest ), // Templated
		       .reg_pipe6_map8_dt_source(reg_pipe6_map8_dt_source ), // Templated
		       .reg_pipe6_map8_vc_dest(reg_pipe6_map8_vc_dest ), // Templated
		       .reg_pipe6_map8_vc_source(reg_pipe6_map8_vc_source ), // Templated
		       .reg_pipe6_map9_aggr_id(reg_pipe6_map9_aggr_id[3:0]),
		       .reg_pipe6_map9_dt_dest(reg_pipe6_map9_dt_dest ), // Templated
		       .reg_pipe6_map9_dt_source(reg_pipe6_map9_dt_source ), // Templated
		       .reg_pipe6_map9_vc_dest(reg_pipe6_map9_vc_dest ), // Templated
		       .reg_pipe6_map9_vc_source(reg_pipe6_map9_vc_source ), // Templated
		       .reg_pipe6_map_en(reg_pipe6_map_en),	 // Templated
		       .reg_pipe6_wr_mode(reg_pipe6_wr_mode[1:0]),
		       .reg_pipe7_drop_ls_le_pkt(reg_pipe7_drop_ls_le_pkt),
		       .reg_pipe7_map0_aggr_id(reg_pipe7_map0_aggr_id[3:0]),
		       .reg_pipe7_map0_dt_dest(reg_pipe7_map0_dt_dest ), // Templated
		       .reg_pipe7_map0_dt_source(reg_pipe7_map0_dt_source ), // Templated
		       .reg_pipe7_map0_vc_dest(reg_pipe7_map0_vc_dest ), // Templated
		       .reg_pipe7_map0_vc_source(reg_pipe7_map0_vc_source ), // Templated
		       .reg_pipe7_map10_aggr_id(reg_pipe7_map10_aggr_id[3:0]),
		       .reg_pipe7_map10_dt_dest(reg_pipe7_map10_dt_dest), // Templated
		       .reg_pipe7_map10_dt_source(reg_pipe7_map10_dt_source), // Templated
		       .reg_pipe7_map10_vc_dest(reg_pipe7_map10_vc_dest), // Templated
		       .reg_pipe7_map10_vc_source(reg_pipe7_map10_vc_source), // Templated
		       .reg_pipe7_map11_aggr_id(reg_pipe7_map11_aggr_id[3:0]),
		       .reg_pipe7_map11_dt_dest(reg_pipe7_map11_dt_dest), // Templated
		       .reg_pipe7_map11_dt_source(reg_pipe7_map11_dt_source), // Templated
		       .reg_pipe7_map11_vc_dest(reg_pipe7_map11_vc_dest), // Templated
		       .reg_pipe7_map11_vc_source(reg_pipe7_map11_vc_source), // Templated
		       .reg_pipe7_map12_aggr_id(reg_pipe7_map12_aggr_id[3:0]),
		       .reg_pipe7_map12_dt_dest(reg_pipe7_map12_dt_dest), // Templated
		       .reg_pipe7_map12_dt_source(reg_pipe7_map12_dt_source), // Templated
		       .reg_pipe7_map12_vc_dest(reg_pipe7_map12_vc_dest), // Templated
		       .reg_pipe7_map12_vc_source(reg_pipe7_map12_vc_source), // Templated
		       .reg_pipe7_map13_aggr_id(reg_pipe7_map13_aggr_id[3:0]),
		       .reg_pipe7_map13_dt_dest(reg_pipe7_map13_dt_dest), // Templated
		       .reg_pipe7_map13_dt_source(reg_pipe7_map13_dt_source), // Templated
		       .reg_pipe7_map13_vc_dest(reg_pipe7_map13_vc_dest), // Templated
		       .reg_pipe7_map13_vc_source(reg_pipe7_map13_vc_source), // Templated
		       .reg_pipe7_map14_aggr_id(reg_pipe7_map14_aggr_id[3:0]),
		       .reg_pipe7_map14_dt_dest(reg_pipe7_map14_dt_dest), // Templated
		       .reg_pipe7_map14_dt_source(reg_pipe7_map14_dt_source), // Templated
		       .reg_pipe7_map14_vc_dest(reg_pipe7_map14_vc_dest), // Templated
		       .reg_pipe7_map14_vc_source(reg_pipe7_map14_vc_source), // Templated
		       .reg_pipe7_map15_aggr_id(reg_pipe7_map15_aggr_id[3:0]),
		       .reg_pipe7_map15_dt_dest(reg_pipe7_map15_dt_dest), // Templated
		       .reg_pipe7_map15_dt_source(reg_pipe7_map15_dt_source), // Templated
		       .reg_pipe7_map15_vc_dest(reg_pipe7_map15_vc_dest), // Templated
		       .reg_pipe7_map15_vc_source(reg_pipe7_map15_vc_source), // Templated
		       .reg_pipe7_map1_aggr_id(reg_pipe7_map1_aggr_id[3:0]),
		       .reg_pipe7_map1_dt_dest(reg_pipe7_map1_dt_dest ), // Templated
		       .reg_pipe7_map1_dt_source(reg_pipe7_map1_dt_source ), // Templated
		       .reg_pipe7_map1_vc_dest(reg_pipe7_map1_vc_dest ), // Templated
		       .reg_pipe7_map1_vc_source(reg_pipe7_map1_vc_source ), // Templated
		       .reg_pipe7_map2_aggr_id(reg_pipe7_map2_aggr_id[3:0]),
		       .reg_pipe7_map2_dt_dest(reg_pipe7_map2_dt_dest ), // Templated
		       .reg_pipe7_map2_dt_source(reg_pipe7_map2_dt_source ), // Templated
		       .reg_pipe7_map2_vc_dest(reg_pipe7_map2_vc_dest ), // Templated
		       .reg_pipe7_map2_vc_source(reg_pipe7_map2_vc_source ), // Templated
		       .reg_pipe7_map3_aggr_id(reg_pipe7_map3_aggr_id[3:0]),
		       .reg_pipe7_map3_dt_dest(reg_pipe7_map3_dt_dest ), // Templated
		       .reg_pipe7_map3_dt_source(reg_pipe7_map3_dt_source ), // Templated
		       .reg_pipe7_map3_vc_dest(reg_pipe7_map3_vc_dest ), // Templated
		       .reg_pipe7_map3_vc_source(reg_pipe7_map3_vc_source ), // Templated
		       .reg_pipe7_map4_aggr_id(reg_pipe7_map4_aggr_id[3:0]),
		       .reg_pipe7_map4_dt_dest(reg_pipe7_map4_dt_dest ), // Templated
		       .reg_pipe7_map4_dt_source(reg_pipe7_map4_dt_source ), // Templated
		       .reg_pipe7_map4_vc_dest(reg_pipe7_map4_vc_dest ), // Templated
		       .reg_pipe7_map4_vc_source(reg_pipe7_map4_vc_source ), // Templated
		       .reg_pipe7_map5_aggr_id(reg_pipe7_map5_aggr_id[3:0]),
		       .reg_pipe7_map5_dt_dest(reg_pipe7_map5_dt_dest ), // Templated
		       .reg_pipe7_map5_dt_source(reg_pipe7_map5_dt_source ), // Templated
		       .reg_pipe7_map5_vc_dest(reg_pipe7_map5_vc_dest ), // Templated
		       .reg_pipe7_map5_vc_source(reg_pipe7_map5_vc_source ), // Templated
		       .reg_pipe7_map6_aggr_id(reg_pipe7_map6_aggr_id[3:0]),
		       .reg_pipe7_map6_dt_dest(reg_pipe7_map6_dt_dest ), // Templated
		       .reg_pipe7_map6_dt_source(reg_pipe7_map6_dt_source ), // Templated
		       .reg_pipe7_map6_vc_dest(reg_pipe7_map6_vc_dest ), // Templated
		       .reg_pipe7_map6_vc_source(reg_pipe7_map6_vc_source ), // Templated
		       .reg_pipe7_map7_aggr_id(reg_pipe7_map7_aggr_id[3:0]),
		       .reg_pipe7_map7_dt_dest(reg_pipe7_map7_dt_dest ), // Templated
		       .reg_pipe7_map7_dt_source(reg_pipe7_map7_dt_source ), // Templated
		       .reg_pipe7_map7_vc_dest(reg_pipe7_map7_vc_dest ), // Templated
		       .reg_pipe7_map7_vc_source(reg_pipe7_map7_vc_source ), // Templated
		       .reg_pipe7_map8_aggr_id(reg_pipe7_map8_aggr_id[3:0]),
		       .reg_pipe7_map8_dt_dest(reg_pipe7_map8_dt_dest ), // Templated
		       .reg_pipe7_map8_dt_source(reg_pipe7_map8_dt_source ), // Templated
		       .reg_pipe7_map8_vc_dest(reg_pipe7_map8_vc_dest ), // Templated
		       .reg_pipe7_map8_vc_source(reg_pipe7_map8_vc_source ), // Templated
		       .reg_pipe7_map9_aggr_id(reg_pipe7_map9_aggr_id[3:0]),
		       .reg_pipe7_map9_dt_dest(reg_pipe7_map9_dt_dest ), // Templated
		       .reg_pipe7_map9_dt_source(reg_pipe7_map9_dt_source ), // Templated
		       .reg_pipe7_map9_vc_dest(reg_pipe7_map9_vc_dest ), // Templated
		       .reg_pipe7_map9_vc_source(reg_pipe7_map9_vc_source ), // Templated
		       .reg_pipe7_map_en(reg_pipe7_map_en),	 // Templated
		       .reg_pipe7_wr_mode(reg_pipe7_wr_mode[1:0]),
		       .reg_pipe_fifo_full_clear(reg_pipe_fifo_full_clear[3:0]),
		       .reg_pipe_fifo_full_clear_last_four(reg_pipe_fifo_full_clear_last_four[3:0]),
		       .reg_resv_pkt_match_lp_dt_en_pipe0(reg_resv_pkt_match_lp_dt_en ), // Templated
		       .reg_resv_pkt_match_lp_dt_en_pipe1(reg_resv_pkt_match_lp_dt_en ), // Templated
		       .reg_resv_pkt_match_lp_dt_en_pipe2(reg_resv_pkt_match_lp_dt_en ), // Templated
		       .reg_resv_pkt_match_lp_dt_en_pipe3(reg_resv_pkt_match_lp_dt_en ), // Templated
		       .reg_resv_pkt_match_lp_dt_en_pipe4(reg_resv_pkt_match_lp_dt_en ), // Templated
		       .reg_resv_pkt_match_lp_dt_en_pipe5(reg_resv_pkt_match_lp_dt_en ), // Templated
		       .reg_resv_pkt_match_lp_dt_en_pipe6(reg_resv_pkt_match_lp_dt_en ), // Templated
		       .reg_resv_pkt_match_lp_dt_en_pipe7(reg_resv_pkt_match_lp_dt_en ), // Templated
		       .reg_resv_pkt_match_lp_dt_pipe0(reg_resv_pkt_match_lp_dt    ), // Templated
		       .reg_resv_pkt_match_lp_dt_pipe1(reg_resv_pkt_match_lp_dt    ), // Templated
		       .reg_resv_pkt_match_lp_dt_pipe2(reg_resv_pkt_match_lp_dt    ), // Templated
		       .reg_resv_pkt_match_lp_dt_pipe3(reg_resv_pkt_match_lp_dt    ), // Templated
		       .reg_resv_pkt_match_lp_dt_pipe4(reg_resv_pkt_match_lp_dt    ), // Templated
		       .reg_resv_pkt_match_lp_dt_pipe5(reg_resv_pkt_match_lp_dt    ), // Templated
		       .reg_resv_pkt_match_lp_dt_pipe6(reg_resv_pkt_match_lp_dt    ), // Templated
		       .reg_resv_pkt_match_lp_dt_pipe7(reg_resv_pkt_match_lp_dt    ), // Templated
		       .reg_sch0_frame_sync_auto_change_pipe_wr_mode(reg_sch0_frame_sync_auto_change_pipe_wr_mode),
		       .reg_sch1_frame_sync_auto_change_pipe_wr_mode(reg_sch1_frame_sync_auto_change_pipe_wr_mode),
		       .reg_sch2_frame_sync_auto_change_pipe_wr_mode(reg_sch2_frame_sync_auto_change_pipe_wr_mode),
		       .reg_sch3_frame_sync_auto_change_pipe_wr_mode(reg_sch3_frame_sync_auto_change_pipe_wr_mode),
		       .reg_sch_data_type_align_fail_int_mask0(1'd0), // Templated
		       .reg_sch_data_type_align_fail_int_mask1(1'd0), // Templated
		       .reg_sch_data_type_align_fail_int_mask2(1'd0), // Templated
		       .reg_sch_data_type_align_fail_int_mask3(1'd0), // Templated
		       .reg_send_pkt_match_lp_dt_aggr0(reg_send_pkt_match_lp_dt    ), // Templated
		       .reg_send_pkt_match_lp_dt_aggr1(reg_send_pkt_match_lp_dt    ), // Templated
		       .reg_send_pkt_match_lp_dt_aggr2(reg_send_pkt_match_lp_dt    ), // Templated
		       .reg_send_pkt_match_lp_dt_aggr3(reg_send_pkt_match_lp_dt    ), // Templated
		       .reg_send_pkt_match_lp_dt_en_aggr0(reg_send_pkt_match_lp_dt_en ), // Templated
		       .reg_send_pkt_match_lp_dt_en_aggr1(reg_send_pkt_match_lp_dt_en ), // Templated
		       .reg_send_pkt_match_lp_dt_en_aggr2(reg_send_pkt_match_lp_dt_en ), // Templated
		       .reg_send_pkt_match_lp_dt_en_aggr3(reg_send_pkt_match_lp_dt_en ), // Templated
		       .reg_sram_lcrc_err_oen(reg_sram_lcrc_err_oen[7:0]),
		       .reg_sync_aggr_0_video_mask_latch_reset(reg_sync_aggr_0_video_mask_latch_reset),
		       .reg_sync_aggr_1_video_mask_latch_reset(reg_sync_aggr_1_video_mask_latch_reset),
		       .reg_sync_aggr_2_video_mask_latch_reset(reg_sync_aggr_2_video_mask_latch_reset),
		       .reg_sync_aggr_3_video_mask_latch_reset(reg_sync_aggr_3_video_mask_latch_reset),
		       .reg_sync_aggr_auto_mask_en(reg_sync_aggr_auto_mask_en[3:0]),
		       .reg_sync_aggr_check_framecount_en(reg_sync_aggr_check_framecount_en),
		       .reg_sync_aggr_check_linecount_en(reg_sync_aggr_check_linecount_en),
		       .reg_sync_aggr_force_video_mask(reg_sync_aggr_force_video_mask[3:0]),
		       .reg_sync_aggr_video_mask_restart(reg_sync_aggr_video_mask_restart[3:0]),
		       .reg_sync_aggr_video_status_info_datatype(reg_sync_aggr_video_status_info_datatype[5:0]),
		       .reg_sync_aggr_video_status_info_linecount(reg_sync_aggr_video_status_info_linecount[15:0]),
		       .reg_sync_aggr_video_status_info_vc(reg_sync_aggr_video_status_info_vc[4:0]),
		       .reg_sync_aggr_video_status_info_wordcount(reg_sync_aggr_video_status_info_wordcount[15:0]),
		       .reg_sync_aggr_video_timeout_threshold(reg_sync_aggr_video_timeout_threshold[19:0]),
		       .reg_testbus_hi8bsel_8bmode(reg_testbus_hi8bsel_8bmode),
		       .reg_testbus_sel_hi0(reg_testbus_sel_hi0[5:0]),
		       .reg_testbus_sel_hi1(reg_testbus_sel_hi1[5:0]),
		       .reg_testbus_sel_lo0(reg_testbus_sel_lo0[5:0]),
		       .reg_testbus_sel_lo1(reg_testbus_sel_lo1[5:0]),
		       .reg_testbus_sel_order0(reg_testbus_sel_order0[3:0]),
		       .reg_testbus_sel_order1(reg_testbus_sel_order1[3:0]),
		       .reg_testbus_sel_swap(reg_testbus_sel_swap[15:0]),
		       .reg_vc_selz_h_mep0(reg_vc_selz_h[7:0]),	 // Templated
		       .reg_vc_selz_h_mep1(reg_vc_selz_h[7:0]),	 // Templated
		       .reg_vc_selz_h_mep2(reg_vc_selz_h[7:0]),	 // Templated
		       .reg_vc_selz_h_mep3(reg_vc_selz_h[7:0]),	 // Templated
		       .reg_vc_selz_l_mep0(reg_vc_selz_l[7:0]),	 // Templated
		       .reg_vc_selz_l_mep1(reg_vc_selz_l[7:0]),	 // Templated
		       .reg_vc_selz_l_mep2(reg_vc_selz_l[7:0]),	 // Templated
		       .reg_vc_selz_l_mep3(reg_vc_selz_l[7:0]),	 // Templated
		       .reg_video_data_fwft_fifo_ovf_int_mask0(reg_video_data_fwft_fifo_ovf_int_mask0),
		       .reg_video_data_fwft_fifo_ovf_int_mask1(reg_video_data_fwft_fifo_ovf_int_mask1),
		       .reg_video_data_fwft_fifo_ovf_int_mask2(reg_video_data_fwft_fifo_ovf_int_mask2),
		       .reg_video_data_fwft_fifo_ovf_int_mask3(reg_video_data_fwft_fifo_ovf_int_mask3),
		       .reg_video_data_fwft_fifo_ovf_int_mask4(reg_video_data_fwft_fifo_ovf_int_mask4),
		       .reg_video_data_fwft_fifo_ovf_int_mask5(reg_video_data_fwft_fifo_ovf_int_mask5),
		       .reg_video_data_fwft_fifo_ovf_int_mask6(reg_video_data_fwft_fifo_ovf_int_mask6),
		       .reg_video_data_fwft_fifo_ovf_int_mask7(reg_video_data_fwft_fifo_ovf_int_mask7),
		       .reg_video_fifo_empty_depend_cnt_mux(reg_video_fifo_empty_depend_cnt_mux),
		       .reg_video_pipe_en(reg_video_pipe_en[7:0]),
		       .reg_vprbs_loopback_app_route_lane0(reg_vprbs_loopback), // Templated
		       .reg_vprbs_loopback_app_route_lane1(reg_vprbs_loopback), // Templated
		       .reg_vprbs_loopback_app_route_lane2(reg_vprbs_loopback), // Templated
		       .reg_vprbs_loopback_app_route_lane3(reg_vprbs_loopback), // Templated
		       .reg_vprbs_loopback_app_route_lane4(reg_vprbs_loopback), // Templated
		       .reg_vprbs_loopback_app_route_lane5(reg_vprbs_loopback), // Templated
		       .reg_vprbs_loopback_app_route_lane6(reg_vprbs_loopback), // Templated
		       .reg_vprbs_loopback_app_route_lane7(reg_vprbs_loopback), // Templated
		       .reg_vprbs_rx_chk_en_app_route_lane0(reg_vprbs_rx_chk_en), // Templated
		       .reg_vprbs_rx_chk_en_app_route_lane1(reg_vprbs_rx_chk_en), // Templated
		       .reg_vprbs_rx_chk_en_app_route_lane2(reg_vprbs_rx_chk_en), // Templated
		       .reg_vprbs_rx_chk_en_app_route_lane3(reg_vprbs_rx_chk_en), // Templated
		       .reg_vprbs_rx_chk_en_app_route_lane4(reg_vprbs_rx_chk_en), // Templated
		       .reg_vprbs_rx_chk_en_app_route_lane5(reg_vprbs_rx_chk_en), // Templated
		       .reg_vprbs_rx_chk_en_app_route_lane6(reg_vprbs_rx_chk_en), // Templated
		       .reg_vprbs_rx_chk_en_app_route_lane7(reg_vprbs_rx_chk_en), // Templated
		       .reg_vprbs_rx_err_clear_app_route_lane0(reg_vprbs_rx_err_clear), // Templated
		       .reg_vprbs_rx_err_clear_app_route_lane1(reg_vprbs_rx_err_clear), // Templated
		       .reg_vprbs_rx_err_clear_app_route_lane2(reg_vprbs_rx_err_clear), // Templated
		       .reg_vprbs_rx_err_clear_app_route_lane3(reg_vprbs_rx_err_clear), // Templated
		       .reg_vprbs_rx_err_clear_app_route_lane4(reg_vprbs_rx_err_clear), // Templated
		       .reg_vprbs_rx_err_clear_app_route_lane5(reg_vprbs_rx_err_clear), // Templated
		       .reg_vprbs_rx_err_clear_app_route_lane6(reg_vprbs_rx_err_clear), // Templated
		       .reg_vprbs_rx_err_clear_app_route_lane7(reg_vprbs_rx_err_clear), // Templated
		       .reg_vprbs_rx_load_app_route_lane0(reg_vprbs_rx_load), // Templated
		       .reg_vprbs_rx_load_app_route_lane1(reg_vprbs_rx_load), // Templated
		       .reg_vprbs_rx_load_app_route_lane2(reg_vprbs_rx_load), // Templated
		       .reg_vprbs_rx_load_app_route_lane3(reg_vprbs_rx_load), // Templated
		       .reg_vprbs_rx_load_app_route_lane4(reg_vprbs_rx_load), // Templated
		       .reg_vprbs_rx_load_app_route_lane5(reg_vprbs_rx_load), // Templated
		       .reg_vprbs_rx_load_app_route_lane6(reg_vprbs_rx_load), // Templated
		       .reg_vprbs_rx_load_app_route_lane7(reg_vprbs_rx_load), // Templated
		       .reg_vprbs_rx_lock_continue_app_route_lane0(reg_vprbs_rx_lock_continue), // Templated
		       .reg_vprbs_rx_lock_continue_app_route_lane1(reg_vprbs_rx_lock_continue), // Templated
		       .reg_vprbs_rx_lock_continue_app_route_lane2(reg_vprbs_rx_lock_continue), // Templated
		       .reg_vprbs_rx_lock_continue_app_route_lane3(reg_vprbs_rx_lock_continue), // Templated
		       .reg_vprbs_rx_lock_continue_app_route_lane4(reg_vprbs_rx_lock_continue), // Templated
		       .reg_vprbs_rx_lock_continue_app_route_lane5(reg_vprbs_rx_lock_continue), // Templated
		       .reg_vprbs_rx_lock_continue_app_route_lane6(reg_vprbs_rx_lock_continue), // Templated
		       .reg_vprbs_rx_lock_continue_app_route_lane7(reg_vprbs_rx_lock_continue), // Templated
		       .reg_vprbs_rx_locked_match_cnt_app_route_lane0(reg_vprbs_rx_locked_match_cnt[3:0]), // Templated
		       .reg_vprbs_rx_locked_match_cnt_app_route_lane1(reg_vprbs_rx_locked_match_cnt[3:0]), // Templated
		       .reg_vprbs_rx_locked_match_cnt_app_route_lane2(reg_vprbs_rx_locked_match_cnt[3:0]), // Templated
		       .reg_vprbs_rx_locked_match_cnt_app_route_lane3(reg_vprbs_rx_locked_match_cnt[3:0]), // Templated
		       .reg_vprbs_rx_locked_match_cnt_app_route_lane4(reg_vprbs_rx_locked_match_cnt[3:0]), // Templated
		       .reg_vprbs_rx_locked_match_cnt_app_route_lane5(reg_vprbs_rx_locked_match_cnt[3:0]), // Templated
		       .reg_vprbs_rx_locked_match_cnt_app_route_lane6(reg_vprbs_rx_locked_match_cnt[3:0]), // Templated
		       .reg_vprbs_rx_locked_match_cnt_app_route_lane7(reg_vprbs_rx_locked_match_cnt[3:0]), // Templated
		       .reg_vprbs_rx_mode_app_route_lane0(reg_vprbs_rx_mode[2:0]), // Templated
		       .reg_vprbs_rx_mode_app_route_lane1(reg_vprbs_rx_mode[2:0]), // Templated
		       .reg_vprbs_rx_mode_app_route_lane2(reg_vprbs_rx_mode[2:0]), // Templated
		       .reg_vprbs_rx_mode_app_route_lane3(reg_vprbs_rx_mode[2:0]), // Templated
		       .reg_vprbs_rx_mode_app_route_lane4(reg_vprbs_rx_mode[2:0]), // Templated
		       .reg_vprbs_rx_mode_app_route_lane5(reg_vprbs_rx_mode[2:0]), // Templated
		       .reg_vprbs_rx_mode_app_route_lane6(reg_vprbs_rx_mode[2:0]), // Templated
		       .reg_vprbs_rx_mode_app_route_lane7(reg_vprbs_rx_mode[2:0]), // Templated
		       .reg_vprbs_rx_order_app_route_lane0(reg_vprbs_rx_order), // Templated
		       .reg_vprbs_rx_order_app_route_lane1(reg_vprbs_rx_order), // Templated
		       .reg_vprbs_rx_order_app_route_lane2(reg_vprbs_rx_order), // Templated
		       .reg_vprbs_rx_order_app_route_lane3(reg_vprbs_rx_order), // Templated
		       .reg_vprbs_rx_order_app_route_lane4(reg_vprbs_rx_order), // Templated
		       .reg_vprbs_rx_order_app_route_lane5(reg_vprbs_rx_order), // Templated
		       .reg_vprbs_rx_order_app_route_lane6(reg_vprbs_rx_order), // Templated
		       .reg_vprbs_rx_order_app_route_lane7(reg_vprbs_rx_order), // Templated
		       .reg_vprbs_rx_uncheck_tolerance_app_route_lane0(reg_vprbs_rx_uncheck_tolerance[3:0]), // Templated
		       .reg_vprbs_rx_uncheck_tolerance_app_route_lane1(reg_vprbs_rx_uncheck_tolerance[3:0]), // Templated
		       .reg_vprbs_rx_uncheck_tolerance_app_route_lane2(reg_vprbs_rx_uncheck_tolerance[3:0]), // Templated
		       .reg_vprbs_rx_uncheck_tolerance_app_route_lane3(reg_vprbs_rx_uncheck_tolerance[3:0]), // Templated
		       .reg_vprbs_rx_uncheck_tolerance_app_route_lane4(reg_vprbs_rx_uncheck_tolerance[3:0]), // Templated
		       .reg_vprbs_rx_uncheck_tolerance_app_route_lane5(reg_vprbs_rx_uncheck_tolerance[3:0]), // Templated
		       .reg_vprbs_rx_uncheck_tolerance_app_route_lane6(reg_vprbs_rx_uncheck_tolerance[3:0]), // Templated
		       .reg_vprbs_rx_uncheck_tolerance_app_route_lane7(reg_vprbs_rx_uncheck_tolerance[3:0]), // Templated
		       .reg_vprbs_tx_err_inject_en_app_route_lane0(reg_vprbs_tx_err_inject_en), // Templated
		       .reg_vprbs_tx_err_inject_en_app_route_lane1(reg_vprbs_tx_err_inject_en), // Templated
		       .reg_vprbs_tx_err_inject_en_app_route_lane2(reg_vprbs_tx_err_inject_en), // Templated
		       .reg_vprbs_tx_err_inject_en_app_route_lane3(reg_vprbs_tx_err_inject_en), // Templated
		       .reg_vprbs_tx_err_inject_en_app_route_lane4(reg_vprbs_tx_err_inject_en), // Templated
		       .reg_vprbs_tx_err_inject_en_app_route_lane5(reg_vprbs_tx_err_inject_en), // Templated
		       .reg_vprbs_tx_err_inject_en_app_route_lane6(reg_vprbs_tx_err_inject_en), // Templated
		       .reg_vprbs_tx_err_inject_en_app_route_lane7(reg_vprbs_tx_err_inject_en), // Templated
		       .reg_vprbs_tx_err_inject_intv_num_app_route_lane0(reg_vprbs_tx_err_inject_intv_num[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_num_app_route_lane1(reg_vprbs_tx_err_inject_intv_num[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_num_app_route_lane2(reg_vprbs_tx_err_inject_intv_num[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_num_app_route_lane3(reg_vprbs_tx_err_inject_intv_num[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_num_app_route_lane4(reg_vprbs_tx_err_inject_intv_num[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_num_app_route_lane5(reg_vprbs_tx_err_inject_intv_num[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_num_app_route_lane6(reg_vprbs_tx_err_inject_intv_num[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_num_app_route_lane7(reg_vprbs_tx_err_inject_intv_num[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_time_app_route_lane0(reg_vprbs_tx_err_inject_intv_time[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_time_app_route_lane1(reg_vprbs_tx_err_inject_intv_time[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_time_app_route_lane2(reg_vprbs_tx_err_inject_intv_time[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_time_app_route_lane3(reg_vprbs_tx_err_inject_intv_time[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_time_app_route_lane4(reg_vprbs_tx_err_inject_intv_time[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_time_app_route_lane5(reg_vprbs_tx_err_inject_intv_time[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_time_app_route_lane6(reg_vprbs_tx_err_inject_intv_time[7:0]), // Templated
		       .reg_vprbs_tx_err_inject_intv_time_app_route_lane7(reg_vprbs_tx_err_inject_intv_time[7:0]), // Templated
		       .reg_vprbs_tx_gen_en_app_route_lane0(reg_vprbs_tx_gen_en), // Templated
		       .reg_vprbs_tx_gen_en_app_route_lane1(reg_vprbs_tx_gen_en), // Templated
		       .reg_vprbs_tx_gen_en_app_route_lane2(reg_vprbs_tx_gen_en), // Templated
		       .reg_vprbs_tx_gen_en_app_route_lane3(reg_vprbs_tx_gen_en), // Templated
		       .reg_vprbs_tx_gen_en_app_route_lane4(reg_vprbs_tx_gen_en), // Templated
		       .reg_vprbs_tx_gen_en_app_route_lane5(reg_vprbs_tx_gen_en), // Templated
		       .reg_vprbs_tx_gen_en_app_route_lane6(reg_vprbs_tx_gen_en), // Templated
		       .reg_vprbs_tx_gen_en_app_route_lane7(reg_vprbs_tx_gen_en), // Templated
		       .reg_vprbs_tx_idi_driver_data_type_app_route_lane0(reg_vprbs_tx_idi_driver_data_type[5:0]), // Templated
		       .reg_vprbs_tx_idi_driver_data_type_app_route_lane1(reg_vprbs_tx_idi_driver_data_type[5:0]), // Templated
		       .reg_vprbs_tx_idi_driver_data_type_app_route_lane2(reg_vprbs_tx_idi_driver_data_type[5:0]), // Templated
		       .reg_vprbs_tx_idi_driver_data_type_app_route_lane3(reg_vprbs_tx_idi_driver_data_type[5:0]), // Templated
		       .reg_vprbs_tx_idi_driver_data_type_app_route_lane4(reg_vprbs_tx_idi_driver_data_type[5:0]), // Templated
		       .reg_vprbs_tx_idi_driver_data_type_app_route_lane5(reg_vprbs_tx_idi_driver_data_type[5:0]), // Templated
		       .reg_vprbs_tx_idi_driver_data_type_app_route_lane6(reg_vprbs_tx_idi_driver_data_type[5:0]), // Templated
		       .reg_vprbs_tx_idi_driver_data_type_app_route_lane7(reg_vprbs_tx_idi_driver_data_type[5:0]), // Templated
		       .reg_vprbs_tx_idi_driver_pkt_interval_app_route_lane0(reg_vprbs_tx_idi_driver_pkt_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_pkt_interval_app_route_lane1(reg_vprbs_tx_idi_driver_pkt_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_pkt_interval_app_route_lane2(reg_vprbs_tx_idi_driver_pkt_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_pkt_interval_app_route_lane3(reg_vprbs_tx_idi_driver_pkt_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_pkt_interval_app_route_lane4(reg_vprbs_tx_idi_driver_pkt_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_pkt_interval_app_route_lane5(reg_vprbs_tx_idi_driver_pkt_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_pkt_interval_app_route_lane6(reg_vprbs_tx_idi_driver_pkt_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_pkt_interval_app_route_lane7(reg_vprbs_tx_idi_driver_pkt_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_total_interval_app_route_lane0(reg_vprbs_tx_idi_driver_total_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_total_interval_app_route_lane1(reg_vprbs_tx_idi_driver_total_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_total_interval_app_route_lane2(reg_vprbs_tx_idi_driver_total_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_total_interval_app_route_lane3(reg_vprbs_tx_idi_driver_total_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_total_interval_app_route_lane4(reg_vprbs_tx_idi_driver_total_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_total_interval_app_route_lane5(reg_vprbs_tx_idi_driver_total_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_total_interval_app_route_lane6(reg_vprbs_tx_idi_driver_total_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_total_interval_app_route_lane7(reg_vprbs_tx_idi_driver_total_interval[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_virtual_channel_app_route_lane0(reg_vprbs_tx_idi_driver_virtual_channel[3:0]), // Templated
		       .reg_vprbs_tx_idi_driver_virtual_channel_app_route_lane1(reg_vprbs_tx_idi_driver_virtual_channel[3:0]), // Templated
		       .reg_vprbs_tx_idi_driver_virtual_channel_app_route_lane2(reg_vprbs_tx_idi_driver_virtual_channel[3:0]), // Templated
		       .reg_vprbs_tx_idi_driver_virtual_channel_app_route_lane3(reg_vprbs_tx_idi_driver_virtual_channel[3:0]), // Templated
		       .reg_vprbs_tx_idi_driver_virtual_channel_app_route_lane4(reg_vprbs_tx_idi_driver_virtual_channel[3:0]), // Templated
		       .reg_vprbs_tx_idi_driver_virtual_channel_app_route_lane5(reg_vprbs_tx_idi_driver_virtual_channel[3:0]), // Templated
		       .reg_vprbs_tx_idi_driver_virtual_channel_app_route_lane6(reg_vprbs_tx_idi_driver_virtual_channel[3:0]), // Templated
		       .reg_vprbs_tx_idi_driver_virtual_channel_app_route_lane7(reg_vprbs_tx_idi_driver_virtual_channel[3:0]), // Templated
		       .reg_vprbs_tx_idi_driver_word_count_app_route_lane0(reg_vprbs_tx_idi_driver_word_count[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_word_count_app_route_lane1(reg_vprbs_tx_idi_driver_word_count[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_word_count_app_route_lane2(reg_vprbs_tx_idi_driver_word_count[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_word_count_app_route_lane3(reg_vprbs_tx_idi_driver_word_count[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_word_count_app_route_lane4(reg_vprbs_tx_idi_driver_word_count[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_word_count_app_route_lane5(reg_vprbs_tx_idi_driver_word_count[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_word_count_app_route_lane6(reg_vprbs_tx_idi_driver_word_count[15:0]), // Templated
		       .reg_vprbs_tx_idi_driver_word_count_app_route_lane7(reg_vprbs_tx_idi_driver_word_count[15:0]), // Templated
		       .reg_vprbs_tx_mode_app_route_lane0(reg_vprbs_tx_mode[2:0]), // Templated
		       .reg_vprbs_tx_mode_app_route_lane1(reg_vprbs_tx_mode[2:0]), // Templated
		       .reg_vprbs_tx_mode_app_route_lane2(reg_vprbs_tx_mode[2:0]), // Templated
		       .reg_vprbs_tx_mode_app_route_lane3(reg_vprbs_tx_mode[2:0]), // Templated
		       .reg_vprbs_tx_mode_app_route_lane4(reg_vprbs_tx_mode[2:0]), // Templated
		       .reg_vprbs_tx_mode_app_route_lane5(reg_vprbs_tx_mode[2:0]), // Templated
		       .reg_vprbs_tx_mode_app_route_lane6(reg_vprbs_tx_mode[2:0]), // Templated
		       .reg_vprbs_tx_mode_app_route_lane7(reg_vprbs_tx_mode[2:0]), // Templated
		       .reg_vprbs_tx_order_app_route_lane0(reg_vprbs_tx_order), // Templated
		       .reg_vprbs_tx_order_app_route_lane1(reg_vprbs_tx_order), // Templated
		       .reg_vprbs_tx_order_app_route_lane2(reg_vprbs_tx_order), // Templated
		       .reg_vprbs_tx_order_app_route_lane3(reg_vprbs_tx_order), // Templated
		       .reg_vprbs_tx_order_app_route_lane4(reg_vprbs_tx_order), // Templated
		       .reg_vprbs_tx_order_app_route_lane5(reg_vprbs_tx_order), // Templated
		       .reg_vprbs_tx_order_app_route_lane6(reg_vprbs_tx_order), // Templated
		       .reg_vprbs_tx_order_app_route_lane7(reg_vprbs_tx_order), // Templated
		       .reg_vprbs_tx_pat_reset_app_route_lane0(reg_vprbs_tx_pat_reset), // Templated
		       .reg_vprbs_tx_pat_reset_app_route_lane1(reg_vprbs_tx_pat_reset), // Templated
		       .reg_vprbs_tx_pat_reset_app_route_lane2(reg_vprbs_tx_pat_reset), // Templated
		       .reg_vprbs_tx_pat_reset_app_route_lane3(reg_vprbs_tx_pat_reset), // Templated
		       .reg_vprbs_tx_pat_reset_app_route_lane4(reg_vprbs_tx_pat_reset), // Templated
		       .reg_vprbs_tx_pat_reset_app_route_lane5(reg_vprbs_tx_pat_reset), // Templated
		       .reg_vprbs_tx_pat_reset_app_route_lane6(reg_vprbs_tx_pat_reset), // Templated
		       .reg_vprbs_tx_pat_reset_app_route_lane7(reg_vprbs_tx_pat_reset), // Templated
		       .treed_reg_bank_clk(treed_reg_bank_clk),
		       .treed_reg_bank_clk_reset_n(treed_reg_bank_clk_reset_n),
		       .mep_clk0	(ppi_clk0),		 // Templated
		       .mep_clk1	(ppi_clk1),		 // Templated
		       .mep_clk2	(ppi_clk2),		 // Templated
		       .mep_clk3	(ppi_clk3),		 // Templated
		       .mep_clk_rst_n0	(ppi_clkrstz0),		 // Templated
		       .mep_clk_rst_n1	(ppi_clkrstz1),		 // Templated
		       .mep_clk_rst_n2	(ppi_clkrstz2),		 // Templated
		       .mep_clk_rst_n3	(ppi_clkrstz3),		 // Templated
		       .reg_pipe0_stream_sel(reg_pipe0_stream_sel[1:0]),
		       .reg_pipe1_stream_sel(reg_pipe1_stream_sel[1:0]),
		       .reg_pipe2_stream_sel(reg_pipe2_stream_sel[1:0]),
		       .reg_pipe3_stream_sel(reg_pipe3_stream_sel[1:0]),
		       .reg_pipe4_stream_sel(reg_pipe4_stream_sel[1:0]),
		       .reg_pipe5_stream_sel(reg_pipe5_stream_sel[1:0]),
		       .reg_pipe6_stream_sel(reg_pipe6_stream_sel[1:0]),
		       .reg_pipe7_stream_sel(reg_pipe7_stream_sel[1:0]),
		       .reg_app_sch0	(reg_app_sch0[15:0]),
		       .reg_app_sch1	(reg_app_sch1[15:0]),
		       .reg_app_sch2	(reg_app_sch2[15:0]),
		       .reg_app_sch3	(reg_app_sch3[15:0]),
		       .reg_time_window0(reg_time_window0[16:0]),
		       .reg_time_window1(reg_time_window1[16:0]),
		       .reg_time_window2(reg_time_window2[16:0]),
		       .reg_time_window3(reg_time_window3[16:0]),
		       .reg_time_window4(reg_time_window4[16:0]),
		       .reg_time_window5(reg_time_window5[16:0]),
		       .reg_time_window6(reg_time_window6[16:0]),
		       .reg_time_window7(reg_time_window7[16:0]),
		       .reg_video_loss_en0(reg_video_loss_en0),
		       .reg_video_loss_en1(reg_video_loss_en1),
		       .reg_video_loss_en2(reg_video_loss_en2),
		       .reg_video_loss_en3(reg_video_loss_en3),
		       .reg_video_loss_en4(reg_video_loss_en4),
		       .reg_video_loss_en5(reg_video_loss_en5),
		       .reg_video_loss_en6(reg_video_loss_en6),
		       .reg_video_loss_en7(reg_video_loss_en7),
		       .reg_line_delay_en0(reg_line_delay_en0),
		       .reg_line_delay_en1(reg_line_delay_en1),
		       .reg_line_delay_en2(reg_line_delay_en2),
		       .reg_line_delay_en3(reg_line_delay_en3),
		       .reg_line_delay_en4(reg_line_delay_en4),
		       .reg_line_delay_en5(reg_line_delay_en5),
		       .reg_line_delay_en6(reg_line_delay_en6),
		       .reg_line_delay_en7(reg_line_delay_en7),
		       .reg_app_aggregation_bypass(reg_app_aggregation_bypass),
		       .reg_sch0_fse_filter(reg_sch0_fse_filter),
		       .reg_sch1_fse_filter(reg_sch1_fse_filter),
		       .reg_sch2_fse_filter(reg_sch2_fse_filter),
		       .reg_sch3_fse_filter(reg_sch3_fse_filter),
		       .mep0_virtual_channel(idi_vc_lane0[1:0]), // Templated
		       .mep1_virtual_channel(idi_vc_lane1[1:0]), // Templated
		       .mep2_virtual_channel(idi_vc_lane2[1:0]), // Templated
		       .mep3_virtual_channel(idi_vc_lane3[1:0]), // Templated
		       .mep0_virtual_channel_x(idi_vcx_lane0[1:0]), // Templated
		       .mep1_virtual_channel_x(idi_vcx_lane1[1:0]), // Templated
		       .mep2_virtual_channel_x(idi_vcx_lane2[1:0]), // Templated
		       .mep3_virtual_channel_x(idi_vcx_lane3[1:0])); // Templated
wire[3:0]idi_virtual_channel_lane0;
assign idi_virtual_channel_lane0 = {idi_vc_lane0,idi_vcx_lane0};

/*  as6s_app  AUTO_TEMPLATE (
        .reg_vpg_bk_lines_qst(vpg_bk_lines_qst0[9:0]),
        .reg_vpg_dt_qst    (vpg_dt_qst0[5:0]),
        .reg_vpg_en    (vpg_en0),
        .reg_vpg_frame_num_mode_qst(vpg_frame_num_mode_qst0[0:0]),
        .reg_vpg_hbp_time_qst(vpg_hbp_time_qst0[11:0]),
        .reg_vpg_hline_time_qst(vpg_hline_time_qst0[14:0]),
        .reg_vpg_hsa_time_qst(vpg_hsa_time_qst0[11:0]),
        .reg_vpg_hsync_packet_en_qst(vpg_hsync_packet_en_qst0),
        .reg_vpg_line_num_mode_qst(vpg_line_num_mode_qst0[1:0]),
        .reg_vpg_max_frame_num_qst(vpg_max_frame_num_qst0[15:0]),
        .reg_vpg_mode_qst    (vpg_mode_qst0),
        .reg_vpg_orientation_qst(vpg_orientation_qst0),
        .reg_vpg_pkt_size_qst(vpg_pkt_size_qst0[13:0]),
        .reg_vpg_start_line_num_qst(vpg_start_line_num_qst0[15:0]),
        .reg_vpg_step_line_num_qst(vpg_step_line_num_qst0[15:0]),
        .reg_vpg_vactive_lines_qst(vpg_vactive_lines_qst0[13:0]),
        .reg_vpg_vbp_lines_qst(vpg_vbp_lines_qst0[9:0]),
        .reg_vpg_vc_qst    (vpg_vc_qst0[1:0]),
        .reg_vpg_vcx_qst    (vpg_vcx_qst0[2:0]),
        .reg_vpg_vfp_lines_qst(vpg_vfp_lines_qst0[9:0]),
        .reg_vpg_vsa_lines_qst(vpg_vsa_lines_qst0[9:0]),
        .app2mep\(.*\)    (),
        .host2app_csi_data                (idi_data_lane0[]),
        .host2app_bytes_en                (idi_byte_en_lane0[]),
        .host2app\(.*\)_data_type            (idi_dt_lane0[]),
        .host2app\(.*\)_virtual_channel        (idi_virtual_channel_lane0[]),
        .host2app\(.*\)    (idi\1_lane@[]),
		.host2app_data_crc	(),
		.reg_rd_vprbs_rx_check_app_lane0(), 
		.reg_rd_vprbs_rx_err_app_lane0(), 
		.reg_rd_vprbs_rx_fail_app_lane0(), 
		.reg_vprbs_\(.*\)_app_lane0(reg_vprbs_\1[]), 
		.reg_rd_dvp_clk_cnt_at_clk_10k(),
		.reg_rd_dvp_pin_square_det_succeed(),

        .reg_resv_pkt_match_lp_dt_en\(.*\)   (reg_resv_pkt_match_lp_dt_en ),
        .reg_resv_pkt_match_lp_dt\(.*\)      (reg_resv_pkt_match_lp_dt    ),
        .reg_clear_resv_pkt_cnt_lp_pf\(.*\)  (reg_clear_resv_pkt_cnt_lp_pf),
        .reg_clear_resv_pkt_cnt_lp_ph\(.*\)  (reg_clear_resv_pkt_cnt_lp_ph),
        .reg_clear_resv_pkt_cnt_sp_fe\(.*\)  (reg_clear_resv_pkt_cnt_sp_fe),
        .reg_clear_resv_pkt_cnt_sp_fs\(.*\)  (reg_clear_resv_pkt_cnt_sp_fs),
        .reg_clear_resv_pkt_cnt_sp_le\(.*\)  (reg_clear_resv_pkt_cnt_sp_le),
        .reg_clear_resv_pkt_cnt_sp_ls\(.*\)  (reg_clear_resv_pkt_cnt_sp_ls),
        .reg_rd_resv_pkt_cnt\(.*\)  (),
		.dvp_pin_d0(pixel_data[0]),
		.dvp_pin_d1(pixel_data[1]),
		.dvp_pin_d2(pixel_data[2]),
		.dvp_pin_d3(pixel_data[3]),
		.dvp_pin_d4(pixel_data[4]),
		.dvp_pin_d5(pixel_data[5]),
		.dvp_pin_d6(pixel_data[6]),
		.dvp_pin_d7(pixel_data[7]),
		.dvp_pin_d8(pixel_data[8]),
		.dvp_pin_d9(pixel_data[9]),
		.dvp_pin_d10(pixel_data[10]),
		.dvp_pin_d11(pixel_data[11]),
		.dvp_pin_d12(pixel_data[12]),
		.dvp_pin_d13(pixel_data[13]),
		.dvp_pin_vs(vsync),
		.dvp_pin_hs(hsync),
		.app2mep_csi_data	(as6s_csi_data[]),
		.app2mep_bytes_en	(as6s_csi_bytes_en[]),
		.app2mep_header_en	(as6s_csi_header_en),
		.app2mep_data_en	(as6s_csi_data_en),
		.app2mep_data_type	(as6s_csi_data_type[]),
		.reg_vpg_data_force_en(1'd0),
		.reg_vpg_data_force_value(1'd0),
        .\(.*\)        (\1[]),
)*/
as6s_app u0_as6s_app(/*autoinst*/
		     // Outputs
		     .reg_rd_dvp_clk_cnt_at_clk_10k(),		 // Templated
		     .reg_rd_dvp_pin_square_det_succeed(),	 // Templated
		     .reg_rd_resv_pkt_cnt_lp_pf_lane0(),	 // Templated
		     .reg_rd_resv_pkt_cnt_lp_ph_lane0(),	 // Templated
		     .reg_rd_resv_pkt_cnt_sp_fe_lane0(),	 // Templated
		     .reg_rd_resv_pkt_cnt_sp_fs_lane0(),	 // Templated
		     .reg_rd_resv_pkt_cnt_sp_le_lane0(),	 // Templated
		     .reg_rd_resv_pkt_cnt_sp_ls_lane0(),	 // Templated
		     .reg_rd_vprbs_rx_check_app_lane0(),	 // Templated
		     .reg_rd_vprbs_rx_err_app_lane0(),		 // Templated
		     .reg_rd_vprbs_rx_fail_app_lane0(),		 // Templated
		     .app2mep_csi_data	(as6s_csi_data[(`MEP_CSI2_HOST_IDI_CSIDATA_SIZE-1):0]), // Templated
		     .app2mep_bytes_en	(as6s_csi_bytes_en[(`MEP_CSI2_HOST_BYTES_EN_SIZE-1):0]), // Templated
		     .app2mep_header_en	(as6s_csi_header_en),	 // Templated
		     .app2mep_data_en	(as6s_csi_data_en),	 // Templated
		     .app2mep_data_type	(as6s_csi_data_type[5:0]), // Templated
		     .app2mep_virtual_channel(),		 // Templated
		     .app2mep_word_count(),			 // Templated
		     .app2mep_ecc	(),			 // Templated
		     .app2mep_dvalid	(),			 // Templated
		     .app2mep_hvalid	(),			 // Templated
		     .app2mep_vvalid	(),			 // Templated
		     .app2mep_data_crc	(),			 // Templated
		     .reg_dvp_mode_en	(reg_dvp_mode_en),	 // Templated
		     .vprbs_rx_fail_app_int(vprbs_rx_fail_app_int), // Templated
		     // Inputs
		     .clk_10K		(clk_10K),		 // Templated
		     .dvp_pin_d0	(pixel_data[0]),	 // Templated
		     .dvp_pin_d1	(pixel_data[1]),	 // Templated
		     .dvp_pin_d10	(pixel_data[10]),	 // Templated
		     .dvp_pin_d11	(pixel_data[11]),	 // Templated
		     .dvp_pin_d12	(pixel_data[12]),	 // Templated
		     .dvp_pin_d13	(pixel_data[13]),	 // Templated
		     .dvp_pin_d2	(pixel_data[2]),	 // Templated
		     .dvp_pin_d3	(pixel_data[3]),	 // Templated
		     .dvp_pin_d4	(pixel_data[4]),	 // Templated
		     .dvp_pin_d5	(pixel_data[5]),	 // Templated
		     .dvp_pin_d6	(pixel_data[6]),	 // Templated
		     .dvp_pin_d7	(pixel_data[7]),	 // Templated
		     .dvp_pin_d8	(pixel_data[8]),	 // Templated
		     .dvp_pin_d9	(pixel_data[9]),	 // Templated
		     .dvp_pin_hs	(hsync),		 // Templated
		     .dvp_pin_vs	(vsync),		 // Templated
		     .reg_app_vc_turn_over_en(reg_app_vc_turn_over_en), // Templated
		     .reg_app_vc_turn_over_mode(reg_app_vc_turn_over_mode), // Templated
		     .reg_clear_resv_pkt_cnt_lp_pf_lane0(reg_clear_resv_pkt_cnt_lp_pf), // Templated
		     .reg_clear_resv_pkt_cnt_lp_ph_lane0(reg_clear_resv_pkt_cnt_lp_ph), // Templated
		     .reg_clear_resv_pkt_cnt_sp_fe_lane0(reg_clear_resv_pkt_cnt_sp_fe), // Templated
		     .reg_clear_resv_pkt_cnt_sp_fs_lane0(reg_clear_resv_pkt_cnt_sp_fs), // Templated
		     .reg_clear_resv_pkt_cnt_sp_le_lane0(reg_clear_resv_pkt_cnt_sp_le), // Templated
		     .reg_clear_resv_pkt_cnt_sp_ls_lane0(reg_clear_resv_pkt_cnt_sp_ls), // Templated
		     .reg_crossbar_0	(reg_crossbar_0[4:0]),	 // Templated
		     .reg_crossbar_1	(reg_crossbar_1[4:0]),	 // Templated
		     .reg_crossbar_10	(reg_crossbar_10[4:0]),	 // Templated
		     .reg_crossbar_11	(reg_crossbar_11[4:0]),	 // Templated
		     .reg_crossbar_12	(reg_crossbar_12[4:0]),	 // Templated
		     .reg_crossbar_13	(reg_crossbar_13[4:0]),	 // Templated
		     .reg_crossbar_14	(reg_crossbar_14[4:0]),	 // Templated
		     .reg_crossbar_15	(reg_crossbar_15[4:0]),	 // Templated
		     .reg_crossbar_16	(reg_crossbar_16[4:0]),	 // Templated
		     .reg_crossbar_17	(reg_crossbar_17[4:0]),	 // Templated
		     .reg_crossbar_18	(reg_crossbar_18[4:0]),	 // Templated
		     .reg_crossbar_19	(reg_crossbar_19[4:0]),	 // Templated
		     .reg_crossbar_2	(reg_crossbar_2[4:0]),	 // Templated
		     .reg_crossbar_20	(reg_crossbar_20[4:0]),	 // Templated
		     .reg_crossbar_21	(reg_crossbar_21[4:0]),	 // Templated
		     .reg_crossbar_22	(reg_crossbar_22[4:0]),	 // Templated
		     .reg_crossbar_23	(reg_crossbar_23[4:0]),	 // Templated
		     .reg_crossbar_3	(reg_crossbar_3[4:0]),	 // Templated
		     .reg_crossbar_4	(reg_crossbar_4[4:0]),	 // Templated
		     .reg_crossbar_5	(reg_crossbar_5[4:0]),	 // Templated
		     .reg_crossbar_6	(reg_crossbar_6[4:0]),	 // Templated
		     .reg_crossbar_7	(reg_crossbar_7[4:0]),	 // Templated
		     .reg_crossbar_8	(reg_crossbar_8[4:0]),	 // Templated
		     .reg_crossbar_9	(reg_crossbar_9[4:0]),	 // Templated
		     .reg_crossbar_hs	(reg_crossbar_hs[4:0]),	 // Templated
		     .reg_crossbar_vs	(reg_crossbar_vs[4:0]),	 // Templated
		     .reg_dbl_mode	(reg_dbl_mode),		 // Templated
		     .reg_de_cnt	(reg_de_cnt[31:0]),	 // Templated
		     .reg_de_high	(reg_de_high[31:0]),	 // Templated
		     .reg_de_low	(reg_de_low[31:0]),	 // Templated
		     .reg_dvp_clk_frequence_det_en(reg_dvp_clk_frequence_det_en), // Templated
		     .reg_dvp_pin_square_det_en(reg_dvp_pin_square_det_en), // Templated
		     .reg_dvp_trigger_en(reg_dvp_trigger_en),	 // Templated
		     .reg_dvp_vprbs_tx_gen_en(reg_dvp_vprbs_tx_gen_en), // Templated
		     .reg_dvp_vprbs_tx_mode(reg_dvp_vprbs_tx_mode[2:0]), // Templated
		     .reg_dvp_vprbs_tx_order(reg_dvp_vprbs_tx_order), // Templated
		     .reg_dvp_vprbs_tx_vs_interval(reg_dvp_vprbs_tx_vs_interval[15:0]), // Templated
		     .reg_force_dvp_data_type(reg_force_dvp_data_type[5:0]), // Templated
		     .reg_force_dvp_virtual_channel(reg_force_dvp_virtual_channel[3:0]), // Templated
		     .reg_force_dvp_word_count(reg_force_dvp_word_count[15:0]), // Templated
		     .reg_force_dvp_word_count_en(reg_force_dvp_word_count_en), // Templated
		     .reg_force_mux_0	(reg_force_mux_0),	 // Templated
		     .reg_force_mux_1	(reg_force_mux_1),	 // Templated
		     .reg_force_mux_10	(reg_force_mux_10),	 // Templated
		     .reg_force_mux_11	(reg_force_mux_11),	 // Templated
		     .reg_force_mux_12	(reg_force_mux_12),	 // Templated
		     .reg_force_mux_13	(reg_force_mux_13),	 // Templated
		     .reg_force_mux_14	(reg_force_mux_14),	 // Templated
		     .reg_force_mux_15	(reg_force_mux_15),	 // Templated
		     .reg_force_mux_16	(reg_force_mux_16),	 // Templated
		     .reg_force_mux_17	(reg_force_mux_17),	 // Templated
		     .reg_force_mux_18	(reg_force_mux_18),	 // Templated
		     .reg_force_mux_19	(reg_force_mux_19),	 // Templated
		     .reg_force_mux_2	(reg_force_mux_2),	 // Templated
		     .reg_force_mux_20	(reg_force_mux_20),	 // Templated
		     .reg_force_mux_21	(reg_force_mux_21),	 // Templated
		     .reg_force_mux_22	(reg_force_mux_22),	 // Templated
		     .reg_force_mux_23	(reg_force_mux_23),	 // Templated
		     .reg_force_mux_3	(reg_force_mux_3),	 // Templated
		     .reg_force_mux_4	(reg_force_mux_4),	 // Templated
		     .reg_force_mux_5	(reg_force_mux_5),	 // Templated
		     .reg_force_mux_6	(reg_force_mux_6),	 // Templated
		     .reg_force_mux_7	(reg_force_mux_7),	 // Templated
		     .reg_force_mux_8	(reg_force_mux_8),	 // Templated
		     .reg_force_mux_9	(reg_force_mux_9),	 // Templated
		     .reg_force_mux_hs	(reg_force_mux_hs),	 // Templated
		     .reg_force_mux_vs	(reg_force_mux_vs),	 // Templated
		     .reg_hs2de_dly	(reg_hs2de_dly[31:0]),	 // Templated
		     .reg_invert_mux_0	(reg_invert_mux_0),	 // Templated
		     .reg_invert_mux_1	(reg_invert_mux_1),	 // Templated
		     .reg_invert_mux_10	(reg_invert_mux_10),	 // Templated
		     .reg_invert_mux_11	(reg_invert_mux_11),	 // Templated
		     .reg_invert_mux_12	(reg_invert_mux_12),	 // Templated
		     .reg_invert_mux_13	(reg_invert_mux_13),	 // Templated
		     .reg_invert_mux_14	(reg_invert_mux_14),	 // Templated
		     .reg_invert_mux_15	(reg_invert_mux_15),	 // Templated
		     .reg_invert_mux_16	(reg_invert_mux_16),	 // Templated
		     .reg_invert_mux_17	(reg_invert_mux_17),	 // Templated
		     .reg_invert_mux_18	(reg_invert_mux_18),	 // Templated
		     .reg_invert_mux_19	(reg_invert_mux_19),	 // Templated
		     .reg_invert_mux_2	(reg_invert_mux_2),	 // Templated
		     .reg_invert_mux_20	(reg_invert_mux_20),	 // Templated
		     .reg_invert_mux_21	(reg_invert_mux_21),	 // Templated
		     .reg_invert_mux_22	(reg_invert_mux_22),	 // Templated
		     .reg_invert_mux_23	(reg_invert_mux_23),	 // Templated
		     .reg_invert_mux_3	(reg_invert_mux_3),	 // Templated
		     .reg_invert_mux_4	(reg_invert_mux_4),	 // Templated
		     .reg_invert_mux_5	(reg_invert_mux_5),	 // Templated
		     .reg_invert_mux_6	(reg_invert_mux_6),	 // Templated
		     .reg_invert_mux_7	(reg_invert_mux_7),	 // Templated
		     .reg_invert_mux_8	(reg_invert_mux_8),	 // Templated
		     .reg_invert_mux_9	(reg_invert_mux_9),	 // Templated
		     .reg_invert_mux_hs	(reg_invert_mux_hs),	 // Templated
		     .reg_invert_mux_vs	(reg_invert_mux_vs),	 // Templated
		     .reg_resv_pkt_match_lp_dt_en_lane0(reg_resv_pkt_match_lp_dt_en ), // Templated
		     .reg_resv_pkt_match_lp_dt_lane0(reg_resv_pkt_match_lp_dt    ), // Templated
		     .reg_vpg_bk_lines_qst(vpg_bk_lines_qst0[9:0]), // Templated
		     .reg_vpg_data_force_en(1'd0),		 // Templated
		     .reg_vpg_data_force_value(1'd0),		 // Templated
		     .reg_vpg_dt_qst	(vpg_dt_qst0[5:0]),	 // Templated
		     .reg_vpg_en	(vpg_en0),		 // Templated
		     .reg_vpg_frame_num_mode_qst(vpg_frame_num_mode_qst0[0:0]), // Templated
		     .reg_vpg_hbp_time_qst(vpg_hbp_time_qst0[11:0]), // Templated
		     .reg_vpg_hline_time_qst(vpg_hline_time_qst0[14:0]), // Templated
		     .reg_vpg_hsa_time_qst(vpg_hsa_time_qst0[11:0]), // Templated
		     .reg_vpg_hsync_packet_en_qst(vpg_hsync_packet_en_qst0), // Templated
		     .reg_vpg_line_num_mode_qst(vpg_line_num_mode_qst0[1:0]), // Templated
		     .reg_vpg_max_frame_num_qst(vpg_max_frame_num_qst0[15:0]), // Templated
		     .reg_vpg_mode_qst	(vpg_mode_qst0),	 // Templated
		     .reg_vpg_orientation_qst(vpg_orientation_qst0), // Templated
		     .reg_vpg_pkt_size_qst(vpg_pkt_size_qst0[13:0]), // Templated
		     .reg_vpg_start_line_num_qst(vpg_start_line_num_qst0[15:0]), // Templated
		     .reg_vpg_step_line_num_qst(vpg_step_line_num_qst0[15:0]), // Templated
		     .reg_vpg_vactive_lines_qst(vpg_vactive_lines_qst0[13:0]), // Templated
		     .reg_vpg_vbp_lines_qst(vpg_vbp_lines_qst0[9:0]), // Templated
		     .reg_vpg_vc_qst	(vpg_vc_qst0[1:0]),	 // Templated
		     .reg_vpg_vcx_qst	(vpg_vcx_qst0[2:0]),	 // Templated
		     .reg_vpg_vfp_lines_qst(vpg_vfp_lines_qst0[9:0]), // Templated
		     .reg_vpg_vsa_lines_qst(vpg_vsa_lines_qst0[9:0]), // Templated
		     .reg_vprbs_loopback_app_lane0(reg_vprbs_loopback), // Templated
		     .reg_vprbs_rx_chk_en_app_lane0(reg_vprbs_rx_chk_en), // Templated
		     .reg_vprbs_rx_err_clear_app_lane0(reg_vprbs_rx_err_clear), // Templated
		     .reg_vprbs_rx_load_app_lane0(reg_vprbs_rx_load), // Templated
		     .reg_vprbs_rx_lock_continue_app_lane0(reg_vprbs_rx_lock_continue), // Templated
		     .reg_vprbs_rx_locked_match_cnt_app_lane0(reg_vprbs_rx_locked_match_cnt[3:0]), // Templated
		     .reg_vprbs_rx_mode_app_lane0(reg_vprbs_rx_mode[2:0]), // Templated
		     .reg_vprbs_rx_order_app_lane0(reg_vprbs_rx_order), // Templated
		     .reg_vprbs_rx_uncheck_tolerance_app_lane0(reg_vprbs_rx_uncheck_tolerance[3:0]), // Templated
		     .reg_vprbs_tx_err_inject_en_app_lane0(reg_vprbs_tx_err_inject_en), // Templated
		     .reg_vprbs_tx_err_inject_intv_num_app_lane0(reg_vprbs_tx_err_inject_intv_num[7:0]), // Templated
		     .reg_vprbs_tx_err_inject_intv_time_app_lane0(reg_vprbs_tx_err_inject_intv_time[7:0]), // Templated
		     .reg_vprbs_tx_gen_en_app_lane0(reg_vprbs_tx_gen_en), // Templated
		     .reg_vprbs_tx_idi_driver_data_type_app_lane0(reg_vprbs_tx_idi_driver_data_type[5:0]), // Templated
		     .reg_vprbs_tx_idi_driver_pkt_interval_app_lane0(reg_vprbs_tx_idi_driver_pkt_interval[15:0]), // Templated
		     .reg_vprbs_tx_idi_driver_total_interval_app_lane0(reg_vprbs_tx_idi_driver_total_interval[15:0]), // Templated
		     .reg_vprbs_tx_idi_driver_virtual_channel_app_lane0(reg_vprbs_tx_idi_driver_virtual_channel[3:0]), // Templated
		     .reg_vprbs_tx_idi_driver_word_count_app_lane0(reg_vprbs_tx_idi_driver_word_count[15:0]), // Templated
		     .reg_vprbs_tx_mode_app_lane0(reg_vprbs_tx_mode[2:0]), // Templated
		     .reg_vprbs_tx_order_app_lane0(reg_vprbs_tx_order), // Templated
		     .reg_vprbs_tx_pat_reset_app_lane0(reg_vprbs_tx_pat_reset), // Templated
		     .reg_vs2de_dly	(reg_vs2de_dly[31:0]),	 // Templated
		     .reg_vs2de_trigger_en(reg_vs2de_trigger_en), // Templated
		     .reg_vs2fe_dly	(reg_vs2fe_dly[31:0]),	 // Templated
		     .reg_vs2fs_dly	(reg_vs2fs_dly[31:0]),	 // Templated
		     .reg_yuyv_mode_en	(reg_yuyv_mode_en),	 // Templated
		     .treed_reg_bank_clk(treed_reg_bank_clk),	 // Templated
		     .treed_reg_bank_clk_reset_n(treed_reg_bank_clk_reset_n), // Templated
		     .app_clk_data	(app_clk_data),		 // Templated
		     .app_clk_rst_n	(app_clk_rst_n),	 // Templated
		     .host2app_csi_data	(idi_data_lane0[(`MEP_CSI2_HOST_IDI_CSIDATA_SIZE-1):0]), // Templated
		     .host2app_bytes_en	(idi_byte_en_lane0[(`MEP_CSI2_HOST_BYTES_EN_SIZE-1):0]), // Templated
		     .host2app_header_en(idi_header_en_lane0),	 // Templated
		     .host2app_data_en	(idi_data_en_lane0),	 // Templated
		     .host2app_data_type(idi_dt_lane0[5:0]),	 // Templated
		     .host2app_virtual_channel(idi_virtual_channel_lane0[(`MEP_CSI2_HOST_VC_WIDTH-1):0]), // Templated
		     .host2app_word_count(idi_word_count_lane0[15:0]), // Templated
		     .host2app_ecc	(idi_ecc_lane0[7:0]),	 // Templated
		     .host2app_dvalid	(idi_dvalid_lane0[(`MEP_CSI2_HOST_N_VIRT_CH-1):0]), // Templated
		     .host2app_hvalid	(idi_hvalid_lane0[(`MEP_CSI2_HOST_N_VIRT_CH-1):0]), // Templated
		     .host2app_vvalid	(idi_vvalid_lane0[(`MEP_CSI2_HOST_N_VIRT_CH-1):0]), // Templated
		     .host2app_data_crc	(),			 // Templated
		     .reg_mem_dt1_selz	(reg_mem_dt1_selz[6:0]), // Templated
		     .reg_mem_dt2_selz	(reg_mem_dt2_selz[6:0]), // Templated
		     .reg_mem_dt7_selz	(reg_mem_dt7_selz[6:0]), // Templated
		     .reg_mem_dt8_selz	(reg_mem_dt8_selz[6:0]), // Templated
		     .reg_mem_dt3_selz	(reg_mem_dt3_selz[7:0]), // Templated
		     .reg_mem_dt4_selz	(reg_mem_dt4_selz[7:0]), // Templated
		     .reg_mem_dt3_selz_en(reg_mem_dt3_selz_en),	 // Templated
		     .reg_mem_dt4_selz_en(reg_mem_dt4_selz_en),	 // Templated
		     .reg_vc_selz_l	(reg_vc_selz_l[7:0]),	 // Templated
		     .reg_vc_selz_h	(reg_vc_selz_h[7:0]),	 // Templated
		     .reg_mipi_host_sel	(reg_mipi_host_sel),	 // Templated
		     .efuse_filedname_valid(efuse_filedname_valid), // Templated
		     .efuse_info_mipi_en(efuse_info_mipi_en),	 // Templated
		     .reg_dvp_mode_en_bank2app(reg_dvp_mode_en_bank2app)); // Templated

/* app_video_prbs_chk   AUTO_TEMPLATE (
    .clk(aggre_clk0),
    .rst_n(aggre_clk_rst_n0),
    .prbs_data_in(idi_prbs_chk_data[127:0]),
    .rx_byte_en(idi_prbs_chk_byte_en[3:0]),
    .rx_data_en(idi_prbs_chk_data_en),
    .rx_header_en(idi_prbs_chk_header_en),
    .rx_data_type(idi_prbs_chk_data_type),
    .reg_vprbs_rx_chk_en	(1'd1),
    .reg_vprbs_rx_mode	(3'd0),
    .reg_vprbs_rx_order	(1'd0),
    .reg_vprbs_rx_load	(1'd1),
	.reg_vprbs_rx_lock_continue(1'd1),
	.reg_vprbs_rx_locked_match_cnt(4'd4),
	.reg_vprbs_rx_uncheck_tolerance(4'd6),
    .reg_vprbs_rx_err_clear(1'd0),
	.reg_rd_vprbs_rx_fail(),
	.reg_rd_vprbs_rx_check(),
	.reg_rd_vprbs_rx_err(),
)*/
app_video_prbs_chk #(
                    .DATA_W(128)
) u_app_video_prbs_chk(/*AUTOINST*/
		       // Outputs
		       .reg_rd_vprbs_rx_check(),		 // Templated
		       .reg_rd_vprbs_rx_fail(),			 // Templated
		       .reg_rd_vprbs_rx_err(),			 // Templated
		       // Inputs
		       .clk		(aggre_clk0),		 // Templated
		       .rst_n		(aggre_clk_rst_n0),	 // Templated
		       .prbs_data_in	(idi_prbs_chk_data[127:0]), // Templated
		       .reg_vprbs_rx_chk_en(1'd1),		 // Templated
		       .reg_vprbs_rx_mode(3'd0),		 // Templated
		       .reg_vprbs_rx_order(1'd0),		 // Templated
		       .reg_vprbs_rx_load(1'd1),		 // Templated
		       .reg_vprbs_rx_lock_continue(1'd1),	 // Templated
		       .reg_vprbs_rx_uncheck_tolerance(4'd6),	 // Templated
		       .reg_vprbs_rx_err_clear(1'd0),		 // Templated
		       .reg_vprbs_rx_locked_match_cnt(4'd4),	 // Templated
		       .rx_byte_en	(idi_prbs_chk_byte_en[3:0]), // Templated
		       .rx_data_en	(idi_prbs_chk_data_en),	 // Templated
		       .rx_header_en	(idi_prbs_chk_header_en), // Templated
		       .rx_data_type	(idi_prbs_chk_data_type)); // Templated

initial begin
    reg_app_wr_idi_data_continue                =   1'd1;
    //as6s_vpg_vc_turn_over
    test_mode                                   =   1'b0;
    reg_app_vc_turn_over_en                     =   1'b1;
    reg_app_vc_turn_over_mode                   =   1'b0;

    reg_last_byte_header_down_mux               =   1'd1; 
    reg_video_fifo_empty_depend_cnt_mux         =   1'd1;
    reg_delete_lp_depend_on_wc_mux              =   1'd1;

    reg_clear_app_full_cnt_async_fifo_pipe0     =   1'd0;
    reg_clear_app_full_cnt_sync_fifo_pipe0      =   1'd0;
    reg_time_window0                            =   17'b0_0000_0000_0011_0010  ;
    reg_video_loss_en0                          =   1'b1                       ;
    reg_line_delay_en0                          =   1'd1                       ;
    reg_clear_app_full_cnt_async_fifo_pipe1     =   1'd0;
    reg_clear_app_full_cnt_sync_fifo_pipe1      =   1'd0;
    reg_time_window1                            =   17'b0_0000_0000_0011_0010  ;
    reg_video_loss_en1                          =   1'b1                       ;
    reg_line_delay_en1                          =   1'd1                       ;
    reg_clear_app_full_cnt_async_fifo_pipe2     =   1'd0;
    reg_clear_app_full_cnt_sync_fifo_pipe2      =   1'd0;
    reg_time_window2                            =   17'b0_0000_0000_0011_0010  ;
    reg_video_loss_en2                          =   1'b1                       ;
    reg_line_delay_en2                          =   1'd1                       ;
    reg_clear_app_full_cnt_async_fifo_pipe3     =   1'd0;
    reg_clear_app_full_cnt_sync_fifo_pipe3      =   1'd0;
    reg_time_window3                            =   17'b0_0000_0000_0011_0010  ;
    reg_video_loss_en3                          =   1'b1                       ;
    reg_line_delay_en3                          =   1'd1                       ;
    reg_clear_app_full_cnt_async_fifo_pipe4     =   1'd0;
    reg_clear_app_full_cnt_sync_fifo_pipe4      =   1'd0;
    reg_time_window4                            =   17'b0_0000_0000_0011_0010  ;
    reg_video_loss_en4                          =   1'b1                       ;
    reg_line_delay_en4                          =   1'd1                       ;
    reg_clear_app_full_cnt_async_fifo_pipe5     =   1'd0;
    reg_clear_app_full_cnt_sync_fifo_pipe5      =   1'd0;
    reg_time_window5                            =   17'b0_0000_0000_0011_0010  ;
    reg_video_loss_en5                          =   1'b1                       ;
    reg_line_delay_en5                          =   1'd1                       ;
    reg_clear_app_full_cnt_async_fifo_pipe6     =   1'd0;
    reg_clear_app_full_cnt_sync_fifo_pipe6      =   1'd0;
    reg_time_window6                            =   17'b0_0000_0000_0011_0010  ;
    reg_video_loss_en6                          =   1'b1                       ;
    reg_line_delay_en6                          =   1'd1                       ;
    reg_clear_app_full_cnt_async_fifo_pipe7     =   1'd0;
    reg_clear_app_full_cnt_sync_fifo_pipe7      =   1'd0;
    reg_time_window7                            =   17'b0_0000_0000_0011_0010  ;
    reg_video_loss_en7                          =   1'b1                       ;
    reg_line_delay_en7                          =   1'd1                       ;

    reg_sch0_fse_filter                         =   1'd0                       ;
    reg_sch1_fse_filter                         =   1'd0                       ;
    reg_sch2_fse_filter                         =   1'd0                       ;
    reg_sch3_fse_filter                         =   1'd0                       ;

    reg_drop_mapping_fault_pkt                  =   8'd0                       ;
    reg_pipe0_drop_ls_le_pkt                    =   1'd0                       ;
    reg_pipe1_drop_ls_le_pkt                    =   1'd0                       ;
    reg_pipe2_drop_ls_le_pkt                    =   1'd0                       ;
    reg_pipe3_drop_ls_le_pkt                    =   1'd0                       ;
    reg_pipe4_drop_ls_le_pkt                    =   1'd0                       ;
    reg_pipe5_drop_ls_le_pkt                    =   1'd0                       ;
    reg_pipe6_drop_ls_le_pkt                    =   1'd0                       ;
    reg_pipe7_drop_ls_le_pkt                    =   1'd0                       ;
    //sync aggre
    reg_sch0_frame_sync_auto_change_pipe_wr_mode = 1'd1;
    reg_sch1_frame_sync_auto_change_pipe_wr_mode = 1'd1;
    reg_sch2_frame_sync_auto_change_pipe_wr_mode = 1'd1;
    reg_sch3_frame_sync_auto_change_pipe_wr_mode = 1'd1;
    reg_app_aggregation_bypass    = 1'd0            ;
    gpio2app_sch0_frame_sync_lock = 1'd0            ;
    gpio2app_sch1_frame_sync_lock = 1'd0            ;
    gpio2app_sch2_frame_sync_lock = 1'd0            ;
    gpio2app_sch3_frame_sync_lock = 1'd0            ;
    reg_app_sch0_frame_sync_lock = 1'd1             ;
    reg_app_sch0_frame_sync_lock_force = 1'd1       ;
    reg_app_sch1_frame_sync_lock = 1'd1             ;
    reg_app_sch1_frame_sync_lock_force = 1'd1       ;
    reg_app_sch2_frame_sync_lock = 1'd1             ;
    reg_app_sch2_frame_sync_lock_force = 1'd1       ;
    reg_app_sch3_frame_sync_lock = 1'd1             ;
    reg_app_sch3_frame_sync_lock_force = 1'd1       ;

    //async aggre
    reg_sch0_frame_sync_lock    = 1'd1              ;
    reg_sch1_frame_sync_lock    = 1'd1              ; 
    reg_sch2_frame_sync_lock    = 1'd1              ; 
    reg_sch3_frame_sync_lock    = 1'd1              ; 

    reg_resv_pkt_match_lp_dt_en  = 1'd0;
    reg_send_pkt_match_lp_dt_en  = 1'd0;
    reg_resv_pkt_match_lp_dt     = 6'd0;
    reg_send_pkt_match_lp_dt     = 6'd0;
    reg_clear_send_pkt_cnt_lp_pf = 1'd0;
    reg_clear_send_pkt_cnt_lp_ph = 1'd0;
    reg_clear_send_pkt_cnt_sp_fe = 1'd0;
    reg_clear_send_pkt_cnt_sp_fs = 1'd0;
    reg_clear_send_pkt_cnt_sp_le = 1'd0;
    reg_clear_send_pkt_cnt_sp_ls = 1'd0;
    reg_clear_resv_pkt_cnt_lp_pf = 1'd0;
    reg_clear_resv_pkt_cnt_lp_ph = 1'd0;
    reg_clear_resv_pkt_cnt_sp_fe = 1'd0;
    reg_clear_resv_pkt_cnt_sp_fs = 1'd0;
    reg_clear_resv_pkt_cnt_sp_le = 1'd0;
    reg_clear_resv_pkt_cnt_sp_ls = 1'd0;

    reg_video_pipe_en            = 8'hff;
    #999950

    reg_clear_resv_pkt_cnt_lp_pf = 1'd1 ;
    reg_clear_resv_pkt_cnt_lp_ph = 1'd1 ;
    reg_clear_resv_pkt_cnt_sp_fe = 1'd1 ;
    reg_clear_resv_pkt_cnt_sp_fs = 1'd1 ;
    reg_clear_resv_pkt_cnt_sp_le = 1'd1 ;
    reg_clear_resv_pkt_cnt_sp_ls = 1'd1 ;
    reg_clear_send_pkt_cnt_lp_pf = 1'd1 ;
    reg_clear_send_pkt_cnt_lp_ph = 1'd1 ;
    reg_clear_send_pkt_cnt_sp_fe = 1'd1 ;
    reg_clear_send_pkt_cnt_sp_fs = 1'd1 ;
    reg_clear_send_pkt_cnt_sp_le = 1'd1 ;
    reg_clear_send_pkt_cnt_sp_ls = 1'd1 ;

end

`include "task_app.v"
//`define ASYNC_M1
initial begin
    //test_cfg
    init_reg_vpg0_random_vc10_test();
    init_reg_vpg1_random_vc10_test();
    init_reg_vpg2_random_vc10_test();
    init_reg_vpg3_random_vc10_test();
    turn_over_vc(2'b00);
    init_reg_as6s_app_filter_turn_off();
    //init_reg_as6s_app_dt_24_pixel();
    //init_reg_as6s_app_filter_vc_dt_0_2b_pixel();
    init_reg_pipe_stream_sel(2'd0,2'd1,2'd2,2'd3,2'd0,2'd1,2'd2,2'd3);

    
    `ifndef SRAM_LCRC_EN
    reg_app_pkt_crc_gen_dis      = 1'h0;
    reg_sram_lcrc_err_oen        = 8'hff;
    reg_app_aggr_idi_crc_chk_en  = 4'hf;
    `else
    reg_app_pkt_crc_gen_dis        = 1'h1;
    reg_sram_lcrc_err_oen        = 8'h00;
    reg_app_aggr_idi_crc_chk_en  = 4'h0;
    `endif

    `ifdef CLK_FORCE_1
    clk_force_1();
    `elsif CLK_FORCE_2
    clk_force_2();
    `elsif CLK_FORCE_SAME
    clk_force_same();
    `elsif CLK_FORCE_1_FPGA
    clk_force_1_fpga();
    `elsif CLK_FORCE_2_FPGA
    clk_force_2_fpga();
    `elsif CLK_FORCE_SAME_FPGA
    clk_force_same_fpga();
    `else 
    clk_force_1();
    `endif

    `ifdef ASYNC_M2_4PIPE_CASE1
    init_reg_async_methed2_4pipe_pipe0123sch12();
    turn_over_vc(2'b01);
    `elsif ASYNC_M2_4PIPE_CASE2
    init_reg_async_methed2_4pipe_pipe01sch1_pipe23sch2();
    turn_over_vc(2'b01);
    `elsif ASYNC_M2_8PIPE_CASE1
    init_reg_async_methed2_8pipe_pipe01234567sch01();
    turn_over_vc(2'b01);
    `elsif ASYNC_M1_4PIPE_CASE1
    init_reg_async_methed1_4pipe_pipe01sch0_pipe23sch1();
    `elsif ASYNC_M1_8PIPE_CASE1
    init_reg_async_methed1_8pipe_pipe0145sch0_pipe2367sch1_case1();
    `elsif ASYNC_M1_8PIPE_CASE2
    init_reg_async_methed1_8pipe_pipe0246sch0_pipe1357sch1_case2();

    `elsif CONCAT_ITLV_4PIPE_CASE1
    init_reg_concat_4pipe_pipesch1();
    `elsif CONCAT_ITLV_4PIPE_CASE2
    init_reg_concat_4pipe_pipe03sch1_pipe12sch2();
    `elsif CONCAT_ITLV_4PIPE_CASE3
    init_reg_concat_4pipe_pipesch1_auto_change_pipe_wr_mode();
    `elsif CONCAT_ITLV_3PIPE_CASE1
    init_reg_concat_3pipe_pipesch1();
    `endif
    //header_en_keep_high_long_time();
    //init_reg_aggr_vc_bit(3'b111,3'b101,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000);
    init_reg_aggr_vc_bit(3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000);
    //modify header_en during time
    //mep0_keep_silence_for_a_while();
    ram_ecc_inject_err();

    `ifdef DVP_RAW10_BYTELOC8
    dvp_raw10_byteloc8();
    `elsif DVP_RAW10_BYTELOC7
    dvp_raw10_byteloc7();
    `elsif DVP_RAW10_BYTELOC6
    dvp_raw10_byteloc6();
    `elsif DVP_RAW10_BYTELOC5
    dvp_raw10_byteloc5();
    `elsif DVP_RAW10_BYTELOC4
    dvp_raw10_byteloc4();
    `elsif DVP_RAW10_BYTELOC3
    dvp_raw10_byteloc3();
    `elsif DVP_RAW10_BYTELOC2
    dvp_raw10_byteloc2();
    `elsif DVP_RAW10_BYTELOC1
    dvp_raw10_byteloc1();
    `elsif DVP_RAW8
    dvp_raw8();
    `elsif DVP_RGB565
    dvp_rgb565();
    `elsif DVP_RAW12_BYTELOC8
    dvp_raw12_byteloc8();
    `elsif DVP_RAW12_BYTELOC7
    dvp_raw12_byteloc7();
    `elsif DVP_RAW12_BYTELOC6
    dvp_raw12_byteloc6();
    `elsif DVP_RAW12_BYTELOC5
    dvp_raw12_byteloc5();
    `elsif DVP_RAW12_BYTELOC4
    dvp_raw12_byteloc4();
    `elsif DVP_RAW12_BYTELOC3
    dvp_raw12_byteloc3();
    `elsif DVP_RAW12_BYTELOC2
    dvp_raw12_byteloc2();
    `elsif DVP_RAW12_BYTELOC1
    dvp_raw12_byteloc1();
    `elsif DVP_RGB888_BYTELOC8
    dvp_rgb888_byteloc8();
    `elsif DVP_RGB888_BYTELOC7
    dvp_rgb888_byteloc7();
    `elsif DVP_RGB888_BYTELOC6
    dvp_rgb888_byteloc6();
    `elsif DVP_RGB888_BYTELOC5
    dvp_rgb888_byteloc5();
    `elsif DVP_RGB888_BYTELOC4
    dvp_rgb888_byteloc4();
    `elsif DVP_RGB888_BYTELOC3
    dvp_rgb888_byteloc3();
    `elsif DVP_RGB888_BYTELOC2
    dvp_rgb888_byteloc2();
    `elsif DVP_RGB888_BYTELOC1
    dvp_rgb888_byteloc1();
    `elsif DVP_YUV422_8BIT_UYVY
    dvp_yuv422_8bit_uyuv();
    `elsif DVP_YUV422_8BIT_YUYV
    dvp_yuv422_8bit_yuyv();
    `elsif DVP_YUV422_8BIT_YUYV_HS_TRIGGER
    dvp_yuv422_8bit_yuyv_hs_trigger();
    `elsif DVP_PRBS_RAW8
    dvp_vprbs_raw8();
    `elsif DVP_ATE_TEST
    dvp_ate_test();
    `endif

end

//****idi random driver

`include "./idi_bus_vip/idi_include.v"

initial begin
    $timeformat(-9 , 6, " ns", 10);
end
//****idi random driver
wire [3:0]      fifo_wrclk                                  ;
wire [3:0]      fifo_wrclk_rst_n                            ;
reg  [1:0]      idi_if_drv_virtual_channel_turn_over [3:0]  ;
wire [3:0]      idi_if_drv_header_en_down                   ;
reg  [3:0]      idi_if_drv_header_en_d1                     ;
genvar          i                                           ;

assign    idi_word_count_lane0    =  test_mode ? idi_vpg_word_count_lane0 : idi_if_drv[0].world_count;
assign    idi_byte_en_lane0       =  test_mode ? idi_vpg_byte_en_lane0    : idi_if_drv[0].byte_en;
assign    idi_header_en_lane0     =  test_mode ? idi_vpg_header_en_lane0  : idi_if_drv[0].header_en;
assign    idi_data_en_lane0       =  test_mode ? idi_vpg_data_en_lane0    : idi_if_drv[0].data_en;
assign    idi_data_lane0          =  test_mode ? idi_vpg_data_lane0       : idi_if_drv[0].csi_data;
assign    idi_vc_lane0            =  test_mode ? idi_vpg_vc_lane0         : idi_if_drv_virtual_channel_turn_over[0];
assign    idi_vcx_lane0           =  test_mode ? idi_vpg_vcx_lane0        : idi_if_drv[0].virtual_channel[3:2];
assign    idi_dt_lane0            =  test_mode ? idi_vpg_dt_lane0         : idi_if_drv[0].data_type;
                                                                            
assign    idi_word_count_lane1    =  test_mode ? idi_vpg_word_count_lane1 : idi_if_drv[1].world_count;
assign    idi_byte_en_lane1       =  test_mode ? idi_vpg_byte_en_lane1    : idi_if_drv[1].byte_en;
assign    idi_header_en_lane1     =  test_mode ? idi_vpg_header_en_lane1  : idi_if_drv[1].header_en;
assign    idi_data_en_lane1       =  test_mode ? idi_vpg_data_en_lane1    : idi_if_drv[1].data_en;
assign    idi_data_lane1          =  test_mode ? idi_vpg_data_lane1       : idi_if_drv[1].csi_data;
assign    idi_vc_lane1            =  test_mode ? idi_vpg_vc_lane1         : idi_if_drv_virtual_channel_turn_over[1];
assign    idi_vcx_lane1           =  test_mode ? idi_vpg_vcx_lane1        : idi_if_drv[1].virtual_channel[3:2];
assign    idi_dt_lane1            =  test_mode ? idi_vpg_dt_lane1         : idi_if_drv[1].data_type;
                                                                            
assign    idi_word_count_lane2    =  test_mode ? idi_vpg_word_count_lane2 : idi_if_drv[2].world_count;
assign    idi_byte_en_lane2       =  test_mode ? idi_vpg_byte_en_lane2    : idi_if_drv[2].byte_en;
assign    idi_header_en_lane2     =  test_mode ? idi_vpg_header_en_lane2  : idi_if_drv[2].header_en;
assign    idi_data_en_lane2       =  test_mode ? idi_vpg_data_en_lane2    : idi_if_drv[2].data_en;
assign    idi_data_lane2          =  test_mode ? idi_vpg_data_lane2       : idi_if_drv[2].csi_data;
assign    idi_vc_lane2            =  test_mode ? idi_vpg_vc_lane2         : idi_if_drv_virtual_channel_turn_over[2];
assign    idi_vcx_lane2           =  test_mode ? idi_vpg_vcx_lane2        : idi_if_drv[2].virtual_channel[3:2];
assign    idi_dt_lane2            =  test_mode ? idi_vpg_dt_lane2         : idi_if_drv[2].data_type;
                                                                            
assign    idi_word_count_lane3    =  test_mode ? idi_vpg_word_count_lane3 : idi_if_drv[3].world_count;
assign    idi_byte_en_lane3       =  test_mode ? idi_vpg_byte_en_lane3    : idi_if_drv[3].byte_en;
assign    idi_header_en_lane3     =  test_mode ? idi_vpg_header_en_lane3  : idi_if_drv[3].header_en;
assign    idi_data_en_lane3       =  test_mode ? idi_vpg_data_en_lane3    : idi_if_drv[3].data_en;
assign    idi_data_lane3          =  test_mode ? idi_vpg_data_lane3       : idi_if_drv[3].csi_data;
assign    idi_vc_lane3            =  test_mode ? idi_vpg_vc_lane3         : idi_if_drv_virtual_channel_turn_over[3];
assign    idi_vcx_lane3           =  test_mode ? idi_vpg_vcx_lane3        : idi_if_drv[3].virtual_channel[3:2];
assign    idi_dt_lane3            =  test_mode ? idi_vpg_dt_lane3         : idi_if_drv[3].data_type;
//
//`include "dump.v"


//turn over idi_if_drv vc channel
assign fifo_wrclk       = {fifo_wrclk3,fifo_wrclk2,fifo_wrclk1,fifo_wrclk0};
assign fifo_wrclk_rst_n = {fifo_wrclk_rst_n3,fifo_wrclk_rst_n2,fifo_wrclk_rst_n1,fifo_wrclk_rst_n0};

generate for(i=0;i<=3;i=i+1)begin:idi_if_drv_header_en_bk
    always@(posedge fifo_wrclk[i] or negedge fifo_wrclk_rst_n[i])begin
        if(~fifo_wrclk_rst_n[i])
            idi_if_drv_header_en_d1[i] <= 1'd0;
        else if(idi_if_drv[i].data_type[5:2] != 4'd0)
            idi_if_drv_header_en_d1[i] <= idi_if_drv[i].header_en;
    end

    assign  idi_if_drv_header_en_down[i] = idi_if_drv_header_en_d1[i] & ~idi_if_drv[i].header_en;

    always@(posedge fifo_wrclk[i] or negedge fifo_wrclk_rst_n[i])begin
        if(~fifo_wrclk_rst_n[i])
            idi_if_drv_virtual_channel_turn_over[i] <= 1'd0;
        else if(idi_if_drv_header_en_down[i])
            idi_if_drv_virtual_channel_turn_over[i] <= (idi_if_drv_virtual_channel_turn_over[i] == 2'd2) ? 2'd0 : idi_if_drv_virtual_channel_turn_over[i] + 1'd1;
    end
end
endgenerate


initial begin
   $fsdbDumpfile("app.fsdb");
   $fsdbDumpvars("+all");
   //$fsdbDumpSVA(0,as6d_app_tb,"+fsdbfile=app.fsdb");
   $fsdbDumpMDA(0, as6d_app_tb);
end


initial begin
    `ifdef SHORT_SIM
    #2ms;
    `else
    #4ms;  
    `endif

    $finish;
end 

//***sva check sch pipe fatal

`ifdef ASYNC_M2
bind as6d_app_tb.u_as6d_app.u_as6d_app_aggregator.u0_as6d_app_aggr_lane.u_as6d_app_pipe_sch.u_as6d_app_pipe_sch_fcfs_m2 sch_chk sch_chk_inst0(0,aggre_clk,up_state_aggre_m2,m2_pipe_ack,m2_pipe_line_end);
bind as6d_app_tb.u_as6d_app.u_as6d_app_aggregator.u1_as6d_app_aggr_lane.u_as6d_app_pipe_sch.u_as6d_app_pipe_sch_fcfs_m2 sch_chk sch_chk_inst1(1,aggre_clk,up_state_aggre_m2,m2_pipe_ack,m2_pipe_line_end);
bind as6d_app_tb.u_as6d_app.u_as6d_app_aggregator.u2_as6d_app_aggr_lane.u_as6d_app_pipe_sch.u_as6d_app_pipe_sch_fcfs_m2 sch_chk sch_chk_inst2(2,aggre_clk,up_state_aggre_m2,m2_pipe_ack,m2_pipe_line_end);
bind as6d_app_tb.u_as6d_app.u_as6d_app_aggregator.u3_as6d_app_aggr_lane.u_as6d_app_pipe_sch.u_as6d_app_pipe_sch_fcfs_m2 sch_chk sch_chk_inst3(3,aggre_clk,up_state_aggre_m2,m2_pipe_ack,m2_pipe_line_end);
`elsif ASYNC_M1                                                                            
bind as6d_app_tb.u_as6d_app.u_as6d_app_aggregator.u0_as6d_app_aggr_lane.u_as6d_app_pipe_sch.u_as6d_app_pipe_sch_fcfs_m1 sch_chk sch_chk_inst0(0,aggre_clk,up_state_aggre,ack_aggre_pre,line_end_aggre);
bind as6d_app_tb.u_as6d_app.u_as6d_app_aggregator.u1_as6d_app_aggr_lane.u_as6d_app_pipe_sch.u_as6d_app_pipe_sch_fcfs_m1 sch_chk sch_chk_inst1(1,aggre_clk,up_state_aggre,ack_aggre_pre,line_end_aggre);
bind as6d_app_tb.u_as6d_app.u_as6d_app_aggregator.u2_as6d_app_aggr_lane.u_as6d_app_pipe_sch.u_as6d_app_pipe_sch_fcfs_m1 sch_chk sch_chk_inst2(2,aggre_clk,up_state_aggre,ack_aggre_pre,line_end_aggre);
bind as6d_app_tb.u_as6d_app.u_as6d_app_aggregator.u3_as6d_app_aggr_lane.u_as6d_app_pipe_sch.u_as6d_app_pipe_sch_fcfs_m1 sch_chk sch_chk_inst3(3,aggre_clk,up_state_aggre,ack_aggre_pre,line_end_aggre);
`elsif AS6D_FILTER_DT_26
bind as6d_app_tb.u0_as6s_app filter_check_dt filter_check_dt_inst0(app_clk_data,reg_mem_dt8_selz[6],reg_mem_dt8_selz[5:0],app2mep_header_en,app2mep_data_type[5:0]);
`endif

`ifdef AS6S_DVP
bind as6d_app_tb.u0_as6s_app dvp_data_chk dvp_data_chk_inst(app_clk_data,app_clk_rst_n,app2mep_header_en,app2mep_data_en,app2mep_csi_data[63:0],app2mep_data_type[5:0]);
`endif


`ifdef APP_CRC_CHECK
reg rand_bit;
initial begin
    rand_bit = 0;
    forever @(posedge fifo_wrclk)begin
        rand_bit = ~rand_bit;
        force   as6d_app_tb.u_as6d_app.u_as6d_app_video_pipe.u0_as6d_app_video_pipe_lane.in_csi_data[0] = rand_bit;
    end
end
`endif


endmodule

module sch_chk(sch_sn,clk,sch_cs,ack,line_end);
    input logic [31:0]  sch_sn        ;
    input logic         clk           ;
    input logic [7:0]   sch_cs        ;
    input logic [7:0]   ack           ;
    input logic [7:0]   line_end      ;
    
    property p_pipe0_check_ack;
        @(posedge clk) (ack[0] |-> (sch_cs == 8'b0000_0001));
    endproperty
    property p_pipe1_check_ack;
        @(posedge clk) (ack[1] |-> (sch_cs == 8'b0000_0010));
    endproperty
    property p_pipe2_check_ack;
        @(posedge clk) (ack[2] |-> (sch_cs == 8'b0000_0100));
    endproperty
    property p_pipe3_check_ack;
        @(posedge clk) (ack[3] |-> (sch_cs == 8'b0000_1000));
    endproperty
    property p_pipe4_check_ack;
        @(posedge clk) (ack[4] |-> (sch_cs == 8'b0001_0000));
    endproperty
    property p_pipe5_check_ack;
        @(posedge clk) (ack[5] |-> (sch_cs == 8'b0010_0000));
    endproperty
    property p_pipe6_check_ack;
        @(posedge clk) (ack[6] |-> (sch_cs == 8'b0100_0000));
    endproperty
    property p_pipe7_check_ack;
        @(posedge clk) (ack[7] |-> (sch_cs == 8'b1000_0000));
    endproperty

    property p_pipe0_check_line_end;
        @(posedge clk) (ack[0] & sch_cs[0] |-> ##[1:$] line_end[0]);
    endproperty
    property p_pipe1_check_line_end;
        @(posedge clk) (ack[1] & sch_cs[1] |-> ##[1:$] line_end[1]);
    endproperty                                                  
    property p_pipe2_check_line_end;                             
        @(posedge clk) (ack[2] & sch_cs[2] |-> ##[1:$] line_end[2]);
    endproperty                                                  
    property p_pipe3_check_line_end;                             
        @(posedge clk) (ack[3] & sch_cs[3] |-> ##[1:$] line_end[3]);
    endproperty                                                  
    property p_pipe4_check_line_end;                             
        @(posedge clk) (ack[4] & sch_cs[4] |-> ##[1:$] line_end[4]);
    endproperty                                                  
    property p_pipe5_check_line_end;                             
        @(posedge clk) (ack[5] & sch_cs[5] |-> ##[1:$] line_end[5]);
    endproperty                                                  
    property p_pipe6_check_line_end;                             
        @(posedge clk) (ack[6] & sch_cs[6] |-> ##[1:$] line_end[6]);
    endproperty                                                  
    property p_pipe7_check_line_end;                             
        @(posedge clk) (ack[7] & sch_cs[7] |-> ##[1:$] line_end[7]);
    endproperty

    a_pipe0_check_ack: assert property (p_pipe0_check_ack)
    else
        $fatal("sch function ack is error,pipe0 sch%d",sch_sn);
    a_pipe1_check_ack: assert property (p_pipe1_check_ack)
    else
        $fatal("sch function ack is error,pipe1 sch%d",sch_sn);
    a_pipe2_check_ack: assert property (p_pipe2_check_ack)
    else
        $fatal("sch function ack is error,pipe2 sch%d",sch_sn);
    a_pipe3_check_ack: assert property (p_pipe3_check_ack)
    else
        $fatal("sch function ack is error,pipe3 sch%d",sch_sn);
    a_pipe4_check_ack: assert property (p_pipe4_check_ack)
    else
        $fatal("sch function ack is error,pipe4 sch%d",sch_sn);
    a_pipe5_check_ack: assert property (p_pipe5_check_ack)
    else
        $fatal("sch function ack is error,pipe5 sch%d",sch_sn);
    a_pipe6_check_ack: assert property (p_pipe6_check_ack)
    else
        $fatal("sch function ack is error,pipe6 sch%d",sch_sn);
    a_pipe7_check_ack: assert property (p_pipe7_check_ack)
    else
        $fatal("sch function ack is error,pipe7 sch%d",sch_sn);


    a_pipe0_check_line_end: assert property (p_pipe0_check_line_end)
    else
        $fatal("sch function line_end is error,pipe0 sch%d",sch_sn);
    a_pipe1_check_line_end: assert property (p_pipe1_check_line_end)
    else
        $fatal("sch function line_end is error,pipe1 sch%d",sch_sn);
    a_pipe2_check_line_end: assert property (p_pipe2_check_line_end)
    else
        $fatal("sch function line_end is error,pipe2 sch%d",sch_sn);
    a_pipe3_check_line_end: assert property (p_pipe3_check_line_end)
    else
        $fatal("sch function line_end is error,pipe3 sch%d",sch_sn);
    a_pipe4_check_line_end: assert property (p_pipe4_check_line_end)
    else
        $fatal("sch function line_end is error,pipe4 sch%d",sch_sn);
    a_pipe5_check_line_end: assert property (p_pipe5_check_line_end)
    else
        $fatal("sch function line_end is error,pipe5 sch%d",sch_sn);
    a_pipe6_check_line_end: assert property (p_pipe6_check_line_end)
    else
        $fatal("sch function line_end is error,pipe6 sch%d",sch_sn);
    a_pipe7_check_line_end: assert property (p_pipe7_check_line_end)
    else
        $fatal("sch function line_end is error,pipe7 sch%d",sch_sn);
endmodule

module filter_check_dt(clk,check_en,filter_dt,vld,dt);
    input logic [5:0]  filter_dt ;
    input logic        vld       ; 
    input logic [5:0]  dt        ;
    input logic        check_en  ;
    input logic        clk       ;

    property s_filter_check_dt;
        @(posedge clk) (check_en&(vld&(dt[5:2]!=4'd0))) |-> (dt == filter_dt);
    endproperty

    a_filter_check_dt: assert property (s_filter_check_dt)
    else
        $fatal("as6s filter_check_dt is error,err dt is %d",dt);

endmodule

module  dvp_data_chk(clk,rst_n,idi_header_en,idi_data_en,idi_data,idi_data_type);
    input logic        clk;
    input logic        rst_n;
    input logic        idi_header_en;
    input logic        idi_data_en;
    input logic [63:0] idi_data;
    input logic [5:0]  idi_data_type;

    property p_dvp_raw10_data_chk;
        @(posedge clk)  disable iff(~rst_n) (idi_header_en && idi_data_en && (idi_data_type == 6'h2B)) |-> ((idi_data == 64'h0000_00ff_0000_0000) ||
                                                                                      (idi_data == 64'h0000_0000_0000_ff00) ||
                                                                                      (idi_data == 64'h00ff_0000_0000_ff00) ||
                                                                                      (idi_data == 64'h0000_0000_ff00_0000) ||
                                                                                      (idi_data == 64'h0000_0000_0000_00ff) ||
                                                                                      (idi_data == 64'h0000_ff00_0000_00ff) ||
                                                                                      (idi_data == 64'h0000_0000_00ff_0000) ||
                                                                                      (idi_data == 64'hff00_0000_00ff_0000));
    endproperty

    property p_dvp_raw12_data_chk;
        @(posedge clk)  disable iff(~rst_n) (idi_header_en && idi_data_en && (idi_data_type == 6'h2C)) |-> ((idi_data == 64'h0000_0000_00ff_0000) ||
                                                                                      (idi_data == 64'h0000_ff00_00ff_0000) ||
                                                                                      (idi_data == 64'h0000_0000_0000_00ff) ||
                                                                                      (idi_data == 64'h0000_0000_ff00_00ff) ||
                                                                                      (idi_data == 64'h00ff_0000_ff00_00ff) ||
                                                                                      (idi_data == 64'h0000_0000_0000_ff00) ||
                                                                                      (idi_data == 64'h0000_00ff_0000_ff00) ||
                                                                                      (idi_data == 64'hff00_00ff_0000_ff00));
    endproperty

    property p_dvp_raw8_data_chk;
        @(posedge clk)  disable iff(~rst_n) (idi_header_en && idi_data_en && (idi_data_type == 6'h2A)) |-> ((idi_data == 64'h0000_0000_0000_0001)||
                                                                                                            (idi_data == 64'h0000_0000_0000_0201)||   
                                                                                                            (idi_data == 64'h0000_0000_0003_0201)||   
                                                                                                            (idi_data == 64'h0000_0000_0403_0201)||   
                                                                                                            (idi_data == 64'h0000_0005_0403_0201)||   
                                                                                                            (idi_data == 64'h0000_0605_0403_0201)||   
                                                                                                            (idi_data == 64'h0007_0605_0403_0201)||   
                                                                                                            (idi_data == 64'h0807_0605_0403_0201));
    endproperty

    property p_dvp_rgb565_data_chk;
        @(posedge clk)  disable iff(~rst_n) (idi_header_en && idi_data_en && (idi_data_type == 6'h2D)) |-> ((idi_data == 64'h0000_0000_0000_4949)||
                                                                                                            (idi_data == 64'h0000_0000_4949_4949)||   
                                                                                                            (idi_data == 64'h0000_4949_4949_4949)||   
                                                                                                            (idi_data == 64'h4949_4949_4949_4949));
    endproperty

    property p_dvp_rgb888_data_chk;
        @(posedge clk)  disable iff(~rst_n) (idi_header_en && idi_data_en && (idi_data_type == 6'h24)) |-> ((idi_data == 64'h0203_0102_0301_0203)||
                                                                                                            (idi_data == 64'h0301_0203_0102_0301)||   
                                                                                                            (idi_data == 64'h0102_0301_0203_0102)||   
                                                                                                            (idi_data == 64'h0000_0000_0001_0203)||   
                                                                                                            (idi_data == 64'h0000_0102_0301_0203)||   
                                                                                                            (idi_data == 64'h0000_0000_0000_0001)||   
                                                                                                            (idi_data == 64'h0000_0000_0102_0301)||   
                                                                                                            (idi_data == 64'h0001_0203_0102_0301)||   
                                                                                                            (idi_data == 64'h0000_0000_0000_0102)||   
                                                                                                            (idi_data == 64'h0000_0001_0203_0102));
    endproperty

    property p_dvp_yuv422_8bit_data_chk;
        @(posedge clk)  disable iff(~rst_n) (idi_header_en && idi_data_en && (idi_data_type == 6'h1e)) |-> ((idi_data == 64'h0201_0301_0201_0301)||
                                                                                                            (idi_data == 64'h0201_0301_0000_0000));
    endproperty

    a_dvp_raw10_data_chk: assert property (p_dvp_raw10_data_chk)
    else
        $fatal("as6s dvp chk is error,datatype is raw10,time is %d",$time);
    a_dvp_raw12_data_chk: assert property (p_dvp_raw12_data_chk)
    else
        $fatal("as6s dvp chk is error,datatype is raw12,time is %d",$time);
    a_dvp_raw8_data_chk: assert property (p_dvp_raw8_data_chk)
    else
        $fatal("as6s dvp chk is error,datatype is raw8,time is %d",$time);
    a_dvp_rgb565_data_chk: assert property (p_dvp_rgb565_data_chk)
    else
        $fatal("as6s dvp chk is error,datatype is rgb565,time is %d",$time);
    a_dvp_rgb888_data_chk: assert property (p_dvp_rgb888_data_chk)
    else
        $fatal("as6s dvp chk is error,datatype is rgb888,time is %d",$time);
    a_dvp_yuv422_8bit_data_chk: assert property (p_dvp_yuv422_8bit_data_chk)
    else
        $fatal("as6s dvp chk is error,datatype is yuv422_8bit,time is %d",$time);

endmodule

