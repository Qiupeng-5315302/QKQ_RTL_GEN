
module ecc_137_top

#

(

    parameter DATA_WIDTH = 137,

    parameter PARITY_WIDTH = 9

)

(

    input   [  DATA_WIDTH-1:0]   data_in,

    output  [  DATA_WIDTH-1:0]   data_out,

    input   [   PARITY_WIDTH-1:0]   parity_in,

    output  [   PARITY_WIDTH-1:0]   parity_out,

    input   bypass,

    output  reg [  DATA_WIDTH-1:0]   mask,

    output  sbit_err,

    output  dbit_err

);



wire  [   PARITY_WIDTH-1:0]   syndrome;

reg   [   1:0]              error;



assign parity_out = ecc_encode(data_in);

assign syndrome = parity_in ^ parity_out;

assign data_out = bypass ? data_in : data_in ^ mask;

assign sbit_err = bypass ? 1'b0 : error[0];

assign dbit_err = bypass ? 1'b0 : error[1];





always @(*)

begin

    error = 2'b00;

    case(syndrome)

    9'b000000000 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b00; end

    9'b100000011 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; error = 2'b01; end

    9'b100000101 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; error = 2'b01; end

    9'b100000110 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; error = 2'b01; end

    9'b000000111 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; error = 2'b01; end

    9'b100001001 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; error = 2'b01; end

    9'b100001010 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; error = 2'b01; end

    9'b000001011 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; error = 2'b01; end

    9'b100001100 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; error = 2'b01; end

    9'b000001101 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; error = 2'b01; end

    9'b000001110 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; error = 2'b01; end

    9'b100001111 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; error = 2'b01; end

    9'b100010001 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; error = 2'b01; end

    9'b100010010 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; error = 2'b01; end

    9'b000010011 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; error = 2'b01; end

    9'b100010100 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; error = 2'b01; end

    9'b000010101 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; error = 2'b01; end

    9'b000010110 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; error = 2'b01; end

    9'b100010111 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; error = 2'b01; end

    9'b100011000 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; error = 2'b01; end

    9'b000011001 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; error = 2'b01; end

    9'b000011010 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; error = 2'b01; end

    9'b100011011 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; error = 2'b01; end

    9'b000011100 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; error = 2'b01; end

    9'b100011101 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; error = 2'b01; end

    9'b100011110 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; error = 2'b01; end

    9'b000011111 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; error = 2'b01; end

    9'b100100001 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; error = 2'b01; end

    9'b100100010 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; error = 2'b01; end

    9'b000100011 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; error = 2'b01; end

    9'b100100100 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; error = 2'b01; end

    9'b000100101 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; error = 2'b01; end

    9'b000100110 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; error = 2'b01; end

    9'b100100111 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; error = 2'b01; end

    9'b100101000 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; error = 2'b01; end

    9'b000101001 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; error = 2'b01; end

    9'b000101010 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; error = 2'b01; end

    9'b100101011 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; error = 2'b01; end

    9'b000101100 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; error = 2'b01; end

    9'b100101101 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; error = 2'b01; end

    9'b100101110 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; error = 2'b01; end

    9'b000101111 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; error = 2'b01; end

    9'b100110000 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; error = 2'b01; end

    9'b000110001 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; error = 2'b01; end

    9'b000110010 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; error = 2'b01; end

    9'b100110011 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; error = 2'b01; end

    9'b000110100 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b100110101 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b100110110 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b000110111 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b000111000 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b100111001 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b100111010 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b000111011 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b100111100 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b000111101 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b000111110 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b100111111 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101000001 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101000010 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001000011 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101000100 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001000101 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001000110 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101000111 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101001000 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001001001 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001001010 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101001011 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001001100 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101001101 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101001110 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001001111 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101010000 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001010001 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001010010 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101010011 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001010100 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101010101 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101010110 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001010111 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001011000 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101011001 : begin mask = 137'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101011010 : begin mask = 137'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001011011 : begin mask = 137'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101011100 : begin mask = 137'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001011101 : begin mask = 137'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001011110 : begin mask = 137'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101011111 : begin mask = 137'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101100000 : begin mask = 137'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001100001 : begin mask = 137'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001100010 : begin mask = 137'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101100011 : begin mask = 137'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001100100 : begin mask = 137'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101100101 : begin mask = 137'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101100110 : begin mask = 137'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001100111 : begin mask = 137'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001101000 : begin mask = 137'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101101001 : begin mask = 137'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101101010 : begin mask = 137'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001101011 : begin mask = 137'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101101100 : begin mask = 137'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001101101 : begin mask = 137'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001101110 : begin mask = 137'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101101111 : begin mask = 137'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001110000 : begin mask = 137'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101110001 : begin mask = 137'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101110010 : begin mask = 137'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001110011 : begin mask = 137'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101110100 : begin mask = 137'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001110101 : begin mask = 137'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001110110 : begin mask = 137'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101110111 : begin mask = 137'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101111000 : begin mask = 137'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001111001 : begin mask = 137'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001111010 : begin mask = 137'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101111011 : begin mask = 137'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001111100 : begin mask = 137'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101111101 : begin mask = 137'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b101111110 : begin mask = 137'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001111111 : begin mask = 137'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b110000001 : begin mask = 137'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b110000010 : begin mask = 137'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b010000011 : begin mask = 137'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b110000100 : begin mask = 137'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b010000101 : begin mask = 137'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b010000110 : begin mask = 137'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b110000111 : begin mask = 137'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b110001000 : begin mask = 137'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b010001001 : begin mask = 137'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b010001010 : begin mask = 137'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b110001011 : begin mask = 137'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b010001100 : begin mask = 137'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b110001101 : begin mask = 137'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b110001110 : begin mask = 137'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b010001111 : begin mask = 137'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b110010000 : begin mask = 137'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b010010001 : begin mask = 137'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b100000000 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b010000000 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b001000000 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b000100000 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b000010000 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b000001000 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b000000100 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b000000010 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    9'b000000001 : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b01; end

    default : begin mask = 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; error = 2'b10; end

    endcase

end



function [  PARITY_WIDTH-1:0] ecc_encode;

    input [ DATA_WIDTH-1:0] d;

    reg [ PARITY_WIDTH-1:0] p;

    begin

    p[0] = d[0] + d[1] + d[3] + d[4] + d[6] + d[8] + d[10] + d[11] + d[13] + d[15] + d[17] + d[19] + d[21] + d[23] + d[25] + d[26] + d[28] + d[30] + d[32] + d[34] + d[36] + d[38] + d[40] + d[42] + d[44] + d[46] + d[48] + d[50] + d[52] + d[54] + d[56] + d[57] + d[59] + d[61] + d[63] + d[65] + d[67] + d[69] + d[71] + d[73] + d[75] + d[77] + d[79] + d[81] + d[83] + d[85] + d[87] + d[89] + d[91] + d[93] + d[95] + d[97] + d[99] + d[101] + d[103] + d[105] + d[107] + d[109] + d[111] + d[113] + d[115] + d[117] + d[119] + d[120] + d[122] + d[124] + d[126] + d[128] + d[130] + d[132] + d[134] + d[136] ;

    p[1] = d[0] + d[2] + d[3] + d[5] + d[6] + d[9] + d[10] + d[12] + d[13] + d[16] + d[17] + d[20] + d[21] + d[24] + d[25] + d[27] + d[28] + d[31] + d[32] + d[35] + d[36] + d[39] + d[40] + d[43] + d[44] + d[47] + d[48] + d[51] + d[52] + d[55] + d[56] + d[58] + d[59] + d[62] + d[63] + d[66] + d[67] + d[70] + d[71] + d[74] + d[75] + d[78] + d[79] + d[82] + d[83] + d[86] + d[87] + d[90] + d[91] + d[94] + d[95] + d[98] + d[99] + d[102] + d[103] + d[106] + d[107] + d[110] + d[111] + d[114] + d[115] + d[118] + d[119] + d[121] + d[122] + d[125] + d[126] + d[129] + d[130] + d[133] + d[134] ;

    p[2] = d[1] + d[2] + d[3] + d[7] + d[8] + d[9] + d[10] + d[14] + d[15] + d[16] + d[17] + d[22] + d[23] + d[24] + d[25] + d[29] + d[30] + d[31] + d[32] + d[37] + d[38] + d[39] + d[40] + d[45] + d[46] + d[47] + d[48] + d[53] + d[54] + d[55] + d[56] + d[60] + d[61] + d[62] + d[63] + d[68] + d[69] + d[70] + d[71] + d[76] + d[77] + d[78] + d[79] + d[84] + d[85] + d[86] + d[87] + d[92] + d[93] + d[94] + d[95] + d[100] + d[101] + d[102] + d[103] + d[108] + d[109] + d[110] + d[111] + d[116] + d[117] + d[118] + d[119] + d[123] + d[124] + d[125] + d[126] + d[131] + d[132] + d[133] + d[134] ;

    p[3] = d[4] + d[5] + d[6] + d[7] + d[8] + d[9] + d[10] + d[18] + d[19] + d[20] + d[21] + d[22] + d[23] + d[24] + d[25] + d[33] + d[34] + d[35] + d[36] + d[37] + d[38] + d[39] + d[40] + d[49] + d[50] + d[51] + d[52] + d[53] + d[54] + d[55] + d[56] + d[64] + d[65] + d[66] + d[67] + d[68] + d[69] + d[70] + d[71] + d[80] + d[81] + d[82] + d[83] + d[84] + d[85] + d[86] + d[87] + d[96] + d[97] + d[98] + d[99] + d[100] + d[101] + d[102] + d[103] + d[112] + d[113] + d[114] + d[115] + d[116] + d[117] + d[118] + d[119] + d[127] + d[128] + d[129] + d[130] + d[131] + d[132] + d[133] + d[134] ;

    p[4] = d[11] + d[12] + d[13] + d[14] + d[15] + d[16] + d[17] + d[18] + d[19] + d[20] + d[21] + d[22] + d[23] + d[24] + d[25] + d[41] + d[42] + d[43] + d[44] + d[45] + d[46] + d[47] + d[48] + d[49] + d[50] + d[51] + d[52] + d[53] + d[54] + d[55] + d[56] + d[72] + d[73] + d[74] + d[75] + d[76] + d[77] + d[78] + d[79] + d[80] + d[81] + d[82] + d[83] + d[84] + d[85] + d[86] + d[87] + d[104] + d[105] + d[106] + d[107] + d[108] + d[109] + d[110] + d[111] + d[112] + d[113] + d[114] + d[115] + d[116] + d[117] + d[118] + d[119] + d[135] + d[136] ;

    p[5] = d[26] + d[27] + d[28] + d[29] + d[30] + d[31] + d[32] + d[33] + d[34] + d[35] + d[36] + d[37] + d[38] + d[39] + d[40] + d[41] + d[42] + d[43] + d[44] + d[45] + d[46] + d[47] + d[48] + d[49] + d[50] + d[51] + d[52] + d[53] + d[54] + d[55] + d[56] + d[88] + d[89] + d[90] + d[91] + d[92] + d[93] + d[94] + d[95] + d[96] + d[97] + d[98] + d[99] + d[100] + d[101] + d[102] + d[103] + d[104] + d[105] + d[106] + d[107] + d[108] + d[109] + d[110] + d[111] + d[112] + d[113] + d[114] + d[115] + d[116] + d[117] + d[118] + d[119] ;

    p[6] = d[57] + d[58] + d[59] + d[60] + d[61] + d[62] + d[63] + d[64] + d[65] + d[66] + d[67] + d[68] + d[69] + d[70] + d[71] + d[72] + d[73] + d[74] + d[75] + d[76] + d[77] + d[78] + d[79] + d[80] + d[81] + d[82] + d[83] + d[84] + d[85] + d[86] + d[87] + d[88] + d[89] + d[90] + d[91] + d[92] + d[93] + d[94] + d[95] + d[96] + d[97] + d[98] + d[99] + d[100] + d[101] + d[102] + d[103] + d[104] + d[105] + d[106] + d[107] + d[108] + d[109] + d[110] + d[111] + d[112] + d[113] + d[114] + d[115] + d[116] + d[117] + d[118] + d[119] ;

    p[7] = d[120] + d[121] + d[122] + d[123] + d[124] + d[125] + d[126] + d[127] + d[128] + d[129] + d[130] + d[131] + d[132] + d[133] + d[134] + d[135] + d[136] ;

    p[8] = d[0] + d[1] + d[2] + d[4] + d[5] + d[7] + d[10] + d[11] + d[12] + d[14] + d[17] + d[18] + d[21] + d[23] + d[24] + d[26] + d[27] + d[29] + d[32] + d[33] + d[36] + d[38] + d[39] + d[41] + d[44] + d[46] + d[47] + d[50] + d[51] + d[53] + d[56] + d[57] + d[58] + d[60] + d[63] + d[64] + d[67] + d[69] + d[70] + d[72] + d[75] + d[77] + d[78] + d[81] + d[82] + d[84] + d[87] + d[88] + d[91] + d[93] + d[94] + d[97] + d[98] + d[100] + d[103] + d[105] + d[106] + d[108] + d[111] + d[112] + d[115] + d[117] + d[118] + d[120] + d[121] + d[123] + d[126] + d[127] + d[130] + d[132] + d[133] + d[135] ;

    ecc_encode = p;

    end

endfunction



endmodule

